��      �yellowbrick.regressor.residuals��ResidualsPlot���)��}�(�force_model���	estimator��sklearn.linear_model._base��LinearRegression���)��}�(�fit_intercept���copy_X���n_jobs�N�positive���n_features_in_�K	�coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK	��h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�CHF�j��)Q?ۛ�j��j?^�]��?>�'R?]�9�h?�Dm�0����I��W?��a
�i�B�&:픎?�t�b�rank_�K	�	singular_�hhK ��h��R�(KK	��h!�CH��0�y�@��#�>Zv@ɛ�M^Ri@����3b@MI;��/T@خ:�N@3�I��{C@�W��i'@�a��w�&@�t�b�
intercept_�h�scalar���h!CvӕW��?���R��_sklearn_version��1.3.0�ub�	is_fitted��auto��name�h�_wrapped�h
�_ax��matplotlib.axes._axes��Axes���)��}�(�_stale���stale_callback�N�_axes�h>�figure��matplotlib.figure��Figure���)��}�(h@�hANhChG�
_transform�N�_transformSet���_visible���	_animated���_alpha�N�clipbox�N�	_clippath�N�_clipon���_label�� ��_picker�N�_rasterized���_agg_filter�N�
_mouseover���
_callbacks��matplotlib.cbook��CallbackRegistry���)��}�(�_signals�]��pchanged�a�exception_handler�hX�_exception_printer����	callbacks�}��_cid_gen�K �_func_cid_map�N�_pickled_cids���ub�_remove_method�N�_url�N�_gid�N�_snap�N�_sketch�N�_path_effects�]��_sticky_edges��matplotlib.artist��_XYPair���]�]������
_in_layout���	_suptitle�N�
_supxlabel�N�
_supylabel�N�_align_label_groups�}�(�x�hX�Grouper���)��}��_mapping�}�sb�y�h�)��}�h�}�sbu�
_localaxes�]�(h>h=)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhi�builtins��getattr���hG�delaxes���R�hjNhkNhlNhmNhnhohphs]�]�����hx��	_position��matplotlib.transforms��Bbox���)��}�(�_parents�}����v�h��TransformedBbox���)��}�(h�}����v�h��BboxTransformTo���)��}�(h�}�(���v�h��CompositeGenericTransform���)��}�(�
input_dims�K�output_dims�Kh�}��P�v�h�)��}�(h�Kh�Kh�}�(�P�v�h��BlendedGenericTransform���)��}�(h�}�(��p�h�)��}�(h�Kh�Kh�}��_invalid�K�_shorthand_name�hR�_a�h��_b�h��ScaledTranslation���)��}�(h�}���p�h�sh�K h�hR�	_inverted�N�_t�K G���8�9���_scale_trans�h��Affine2D���)��}�(h�}�(���k�h�)��}�(h�}���k�h�)��}�(h�}�(�оt�h�)��}�(h�}���Lu�h�)��}�(h�}�(�Pr�h�)��}�(h�Kh�Kh�}��P�h�h�)��}�(h�Kh�Kh�}�(�ʙ�h�)��}�(h�}�(��"{�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}���"{�h�sh�K h�hRh�Nh�K G���8�9��h�hό_mtx�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bubub�Ps�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��Ps�h�sh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nubub��5{�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}���5{�h�sh�K h�hRh�Nh�K G���8�9��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bubub�P<{�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��P<{�j	  sh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nubub�м|�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��м|�j  sh�Kh�hRh�Nh�K G��-��-�؆�h�h�h�Nubub�P}�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��P}�j  sh�Kh�hRh�Nh�K G?�-��-�؆�h�h�h�Nubub�J��h��TransformedPath���)��}�(h�}�h�Kh�hR�_path��matplotlib.path��Path���)��}�(�	_vertices�hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�b�_codes�N�_interpolation_steps�K��_simplify_threshold�G?�q�q�֌_should_simplify���	_readonly��ubhIh�_transformed_path�j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ub�_transformed_points�j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P]��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P`��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub� ��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��i�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�)��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        @       @              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub���]�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       @      @              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��+}�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       @      @              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ububuh�Kh�hR�_x�h�_y�hی_affine�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CHŠk�.p@        
�J�\�             xz@9��8��I@                      �?�t�bubub���h�)��}�(h�}�(�P�i�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}��P�i�j�  sh�K h�hRh�Nh�G���8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#�              �?                              �?�t�bubub���|�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}����|�j�  sh�Kh�hRh�Nh�G?��8�9K ��h�h�h�Nubub���|�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}����|�j�  sh�K h�hRh�Nh�G���8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#�              �?                              �?�t�bubub���|�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}����|�j�  sh�Kh�hRh�Nh�G?��8�9K ��h�h�h�Nubub��yz�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}���yz�j�  sh�Kh�hRh�Nh�G��-��-��K ��h�h�h�Nubub�xz�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}��xz�j�  sh�Kh�hRh�Nh�G?�-��-��K ��h�h�h�Nubub��~�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubub���|�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�433333㿔t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Э��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ٿ������ٿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�N��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ɿ������ɿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��yq�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Y�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j;  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j;  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub����j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  jJ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jJ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�bq�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�?433333�?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  jY  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jY  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ububuh�Kh�hRj�  h�j�  h�j�  h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@        ���@;t@����l�o@                      �?�t�bububuh�Kh�hRh�h��TransformWrapper���)��}�(h�}�(�Pcu�h�)��}�(h�}���
�h��BboxTransformFrom���)��}�(h�}��Pr�h�sh�K h�hRh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH��l%��?        �Ԓ.�p�?        �v����?����p�                      �?�t�bub�_boxin�jo  h�hhK ��h��R�(KKK��h!�CH�!��>�?        ��d*R�ֿ        ��tSau�?�S�Ġ��?                      �?�t�bubsh�K h�hR�_bbox�h�)��}�(h�}��Pcu�jo  sh�K h�hR�_points�hhK ��h��R�(KKK��h!�C �Ԓ.�p�?����p俲[8^@�J�Qv��?�t�b�_minpos�hhK ��h��R�(KK��h!�C      �      ��t�b�_ignore���_points_orig�hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjl  j�  hhK ��h��R�(KKK��h!�C �Ԓ.�p�?����p俲[8^@�J�Qv��?�t�bub�P�h�h�uh�K h�hR�_child�h��BlendedAffine2D���)��}�(h�}��Pdu�jl  sh�K h�hRj�  h��IdentityTransform���)��}�(h�}���y�j�  sh�Kh�hRh�Nubj�  j�  )��}�(h�}���y�j�  sh�Kh�hRh�Nubh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bub�	transform�h�j�  j�  ��R��transform_affine�h�j�  j�  ��R��transform_non_affine�h�j�  j�  ��R��transform_path�h�j�  j�  ��R��transform_path_affine�h�j�  j�  ��R��transform_path_non_affine�h�j�  j�  ��R��
get_affine�h�j�  j�  ��R��inverted�h�j�  j�  ��R��
get_matrix�h�j�  j�  ��R�ubh�h�ubsh�Kh�hRh�jt  h�h�ub�ʙ�h���j�  ��Yn�j�  )��}�(h�}�h�Kh�hRj�  j�  )��}�(h�}���Yn�j�  sh�Kh�hRh�Nubj�  h�h�Nh�hhK ��h��R�(KKK��h!�CH      �?                             xz@9��8��I@                      �?�t�bub��s�j�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}���s�j�  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@              �?                              �?�t�bub�P'r�j�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}��P'r�j�  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@              �?                              �?�t�bub�\e�j�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}��\e�j  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH     �@              Y@              �?                              �?�t�bub��|�h�)��}�(h�Kh�Kh�}����|�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����|�j  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���|�j  sh�Kh�hRh�h�)��}�(h�}����|�j*  sh�Kh�hRh�N�_boxout�h�)��}�(h�}���jz�j-  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}����|�j*  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���|�h�)��}�(h�Kh�Kh�}��P}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P}�jR  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjO  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����|�jO  sh�Kh�hRh�h�)��}�(h�}���}�jj  sh�Kh�hRh�Nj0  h�)��}�(h�}���}�jm  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���}�jj  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��}�h�)��}�(h�Kh�Kh�}���}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���}�j�  sh�Kh�hRh�h�)��}�(h�}��}�j�  sh�K h�hRh�Nj0  h�)��}�(h�}��}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��}�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P#}�h�)��}�(h�Kh�Kh�}���#}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���#}�j�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P#}�j�  sh�Kh�hRh�h�)��}�(h�}���"}�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}���!}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���"}�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�'}�h�)��}�(h�Kh�Kh�}��P'}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P'}�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��'}�j  sh�Kh�hRh�h�)��}�(h�}���&}�j9  sh�K h�hRh�Nj0  h�)��}�(h�}���%}�j<  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���&}�j9  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���|�h�)��}�(h�Kh�Kh�}���|�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���|�jf  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjc  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����|�jc  sh�Kh�hRh�h�)��}�(h�}��P�|�j~  sh�Kh�hRh�Nj0  h�)��}�(h�}��P)}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P�|�j~  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�|�h�)��}�(h�Kh�Kh�}��P�|�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�|�j�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�|�j�  sh�Kh�hRh�h�)��}�(h�}���|�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}����|�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���|�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��3{�h�)��}�(h�Kh�Kh�}��P4{�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P4{�j�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���3{�j�  sh�Kh�hRh�h�)��}�(h�}��P�|�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}��P��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P�|�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pjz�h�)��}�(h�Kh�Kh�}��Pfz�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pfz�j#  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj   j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pjz�j   sh�Kh�hRh�h�)��}�(h�}��Prz�j;  sh�Kh�hRh�Nj0  h�)��}�(h�}��zz�j>  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��Prz�j;  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��?y�h�)��}�(h�Kh�Kh�}��P(y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P(y�jb  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj_  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���?y�j_  sh�Kh�hRh�h�)��}�(h�}���y�j�  sh�K h�hRh�Nj0  h�)��}�(h�}��Pz��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���y�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P9y�h�)��}�(h�Kh�Kh�}��P&y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P&y�j�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P9y�j�  sh�Kh�hRh�h�)��}�(h�}��P1y�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}���!y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P1y�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�3y�h�)��}�(h�Kh�Kh�}���y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��3y�j�  sh�Kh�hRh�h�)��}�(h�}���+y�j
  sh�K h�hRh�Nj0  h�)��}�(h�}���&y�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���+y�j
  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��%y�h�)��}�(h�Kh�Kh�}��y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��y�j7  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj4  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���%y�j4  sh�Kh�hRh�h�)��}�(h�}��0y�jO  sh�Kh�hRh�Nj0  h�)��}�(h�}��P5y�jR  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��0y�jO  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�6y�h�)��}�(h�Kh�Kh�}��� y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��� y�jv  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjs  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��6y�js  sh�Kh�hRh�h�)��}�(h�}���4y�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}���?y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���4y�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j�  sh�Kh�hRh�h�)��}�(h�}���y�j�  sh�K h�hRh�Nj0  h�)��}�(h�}��нy�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���y�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��T��h�)��}�(h�Kh�Kh�}��PV��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PV��j   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���T��j�  sh�Kh�hRh�h�)��}�(h�}���U��j  sh�K h�hRh�Nj0  h�)��}�(h�}��PT��j!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���U��j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�в��h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}�(�в��jH  ��i�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�jK  ub�P�|�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�jK  ubuh�K h�hRh�Nh�G        G?�UUUUUU��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?������ @                      �?�t�bubub��i�jN  �P�|�jQ  ���h�)��}�(h�Kh�Kh�}��Sz�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Sz�j^  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj[  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����j[  sh�Kh�hRh�h�)��}�(h�}���f��j|  sh�K h�hRh�Nj0  h�)��}�(h�}��Гy�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���f��j|  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ubuh�Kh�hRh�Nj0  h�h�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@             xz@9��8��I@                      �?�t�bubsh�Kh�hRj�  h�)��}�(h�}��оt�h�sh�K h�hRj�  hhK ��h��R�(KKK��h!�C       �?(\���(�?ffffff�?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIh�j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bub���v�h�uh�Kh�hRh�Nj0  h�h�hhK ��h��R�(KKK��h!�CH      �@        �q�q�@�             0�@�q�q"�                      �?�t�bubsh�K h�hRj�  h�)��}�(h�}����k�h�sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                        @      @�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                        @      @�t�bubhIh�j�  hhK ��h��R�(KKK��h!�C                       �@     0�@�t�bub�PU�h�P+y�h��Py�h���:{�j  ��e�j�  �Ж|�j�  �l�j�  ��{�j�  ��{�j  ��}�j  ��{�j�  �PAz�j�  ��Nq�hƊP
y�h�)��}�(h�}����v�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nub��}z�h�)��}�(h�}����p�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�K h�hRh�Nh�K G���8�9��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bub�Ђp�h�)��}�(h�}��Жp�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nub�Pnz�h�)��}�(h�}���xu�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�)��}�(h�}�(��xu�j  ��u�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}���u�j  sh�K h�hRh�Nh�G?��8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#@              �?                              �?�t�bubub�Oq�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}��Oq�j  sh�Kh�hRh�Nh�G���8�9K ��h�h�h�Nubub�лe�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}��лe�j   sh�K h�hRh�Nh�G?��8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#@              �?                              �?�t�bubub��oz�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}���oz�j-  sh�Kh�hRh�Nh�G��-��-��K ��h�h�h�Nubub�Мy�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}��Мy�j4  sh�Kh�hRh�Nh�G?�-��-��K ��h�h�h�Nubub�P���j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubj8  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubub�����j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�433333㿔t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Pӏ�j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ٿ������ٿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�����j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ɿ������ɿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub���j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�����j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Е��j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub����j  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�?433333�?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ububuh�Kh�hRj�  h�j�  h�j�  h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �8��8V�@        ���@;t@����l�o@                      �?�t�bububh�j  ubsh�Kh�hRh�Nh�G���8�9K ��h�h�h�Nub�yu�j  ��Lz�j  �s�j#  ��Eq�h�)��}�(h�}�(�r�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ub���r�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ub��i�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubuh�K h�hRh�Nh�G        G?�UUUUUU��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?������ @                      �?�t�bub�P�l�h�)��}�(h�}���!t�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G��-��-�؆�h�h�h�Nub��}�h�)��}�(h�}���*}�h�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G?�-��-�؆�h�h�h�Nub��h�j0  �P�y�j7  ��݀�jK  uh�K h�hRh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH{�G�z�?                        {�G�z�?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      Y@                              Y@                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bubub���v�j�  ���p�j�  �Жp�j�  ��!t�j�  ��*}�j�  uh�Kh�hRj�  h�j�  h�j�  h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CHn�d���@        �8��8V�@             xz@9��8��I@                      �?�t�bubub�P�v�j	  uh�Kh�hRh�jk  )��}�(h�}�(���v�h�)��}�(h�}��P�v�js  )��}�(h�}����v�h�sh�K h�hRh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH33333�F@                        �v����?����p�                      �?�t�bubj�  j�  h�hhK ��h��R�(KKK��h!�CH�����?               �        ��tSau�?�S�Ġ��?                      �?�t�bubsh�K h�hRj�  h�)��}�(h�}����v�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C         ����p�33333�F@�J�Qv��?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C         ����p�33333�F@�J�Qv��?�t�bub�P�v�h�uh�K h�hRj�  j�  )��}�(h�}��P�v�j�  sh�K h�hRj�  j�  )��}�(h�}��P�|�j/	  sh�Kh�hRh�Nubj�  j�  )��}�(h�}��P�|�j/	  sh�Kh�hRh�Nubh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�j�  ubj�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�ubh�h�ubsh�Kh�hRh�j	  h�h�ub�P�v�h��P�v�j	  ��1{�j�  )��}�(h�}�h�Kh�hRj�  j�  )��}�(h�}���1{�jS	  sh�Kh�hRh�Nubj�  h�h�Nh�hhK ��h��R�(KKK��h!�CH      �?                             xz@�����?N@                      �?�t�bub��v�j�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}���v�j_	  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �����_�@              �?                              �?�t�bub�dz�j�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}��dz�jk	  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �8��8V�@              �?                              �?�t�bub�P�|�j�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}��P�|�jw	  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �����_�@              �?                              �?�t�bub�r�j�  ���r�j�  ��i�j�  ��y�h�)��}�(h�Kh�Kh�}���l�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���l�j�	  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�	  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���y�j�	  sh�Kh�hRh�h�)��}�(h�}���*{�j�	  sh�Kh�hRh�Nj0  h�)��}�(h�}��]q�j�	  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���*{�j�	  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��.}�h�)��}�(h�Kh�Kh�}���.}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���.}�j�	  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�	  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���.}�j�	  sh�Kh�hRh�h�)��}�(h�}���,}�j�	  sh�Kh�hRh�Nj0  h�)��}�(h�}��P,}�j�	  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���,}�j�	  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��1}�h�)��}�(h�Kh�Kh�}��2}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��2}�j
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���1}�j
  sh�Kh�hRh�h�)��}�(h�}��P1}�j
  sh�Kh�hRh�Nj0  h�)��}�(h�}��P0}�j
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P1}�j
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��5}�h�)��}�(h�Kh�Kh�}���5}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���5}�jC
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj@
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���5}�j@
  sh�Kh�hRh�h�)��}�(h�}��5}�j[
  sh�Kh�hRh�Nj0  h�)��}�(h�}��4}�j^
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��5}�j[
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P9}�h�)��}�(h�Kh�Kh�}���9}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���9}�j�
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P9}�j
  sh�Kh�hRh�h�)��}�(h�}���8}�j�
  sh�Kh�hRh�Nj0  h�)��}�(h�}���7}�j�
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���8}�j�
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�=}�h�)��}�(h�Kh�Kh�}��P=}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P=}�j�
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��=}�j�
  sh�Kh�hRh�h�)��}�(h�}���<}�j�
  sh�Kh�hRh�Nj0  h�)��}�(h�}���;}�j�
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���<}�j�
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��y�h�)��}�(h�Kh�Kh�}��P�y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�y�j   sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���y�j�
  sh�Kh�hRh�h�)��}�(h�}����y�j  sh�Kh�hRh�Nj0  h�)��}�(h�}��P?}�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}����y�j  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���y�h�)��}�(h�Kh�Kh�}��Єy�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Єy�j?  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj<  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����y�j<  sh�Kh�hRh�h�)��}�(h�}���y�jW  sh�Kh�hRh�Nj0  h�)��}�(h�}���y�jZ  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���y�jW  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Фy�h�)��}�(h�Kh�Kh�}���y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���y�j~  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj{  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Фy�j{  sh�Kh�hRh�h�)��}�(h�}����y�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}����y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}����y�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��y�h�)��}�(h�Kh�Kh�}��P�y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���y�j�  sh�Kh�hRh�h�)��}�(h�}����y�j�  sh�K h�hRh�Nj0  h�)��}�(h�}����y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����y�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Ыy�h�)��}�(h�Kh�Kh�}���y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���y�j  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Ыy�j  sh�Kh�hRh�h�)��}�(h�}��P�y�j   sh�Kh�hRh�Nj0  h�)��}�(h�}��P�y�j#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P�y�j   sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���y�h�)��}�(h�Kh�Kh�}��Яy�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Яy�jG  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjD  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����y�jD  sh�Kh�hRh�h�)��}�(h�}���y�je  sh�K h�hRh�Nj0  h�)��}�(h�}���y�jh  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���y�je  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�y�h�)��}�(h�Kh�Kh�}����y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����y�j�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�y�j�  sh�Kh�hRh�h�)��}�(h�}��вy�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}��бy�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��вy�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��y�h�)��}�(h�Kh�Kh�}��P�y�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�y�j�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���y�j�  sh�Kh�hRh�h�)��}�(h�}����y�j�  sh�Kh�hRh�Nj0  h�)��}�(h�}����y�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}����y�j�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j  sh�Kh�hRh�h�)��}�(h�}��P�}�j.  sh�K h�hRh�Nj0  h�)��}�(h�}���_z�j1  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�}�j.  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}���}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���}�j[  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjX  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�jX  sh�Kh�hRh�h�)��}�(h�}����}�jy  sh�K h�hRh�Nj0  h�)��}�(h�}����}�j|  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����}�jy  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j�  sh�Kh�hRh�h�)��}�(h�}���}�j�  sh�K h�hRh�Nj0  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���}�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���}�j�  sh�Kh�hRh�h�)��}�(h�}���}�j  sh�K h�hRh�Nj0  h�)��}�(h�}���}�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���}�j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}���}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���}�j<  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj9  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j9  sh�Kh�hRh�h�)��}�(h�}����}�jZ  sh�K h�hRh�Nj0  h�)��}�(h�}��P�}�j]  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����}�jZ  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}��P�}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j�  sh�Kh�hRh�h�)��}�(h�}����}�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����}�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j�  sh�Kh�hRh�h�)��}�(h�}��P�}�j�  sh�K h�hRh�Nj0  h�)��}�(h�}��P�}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�}�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��}�h�)��}�(h�Kh�Kh�}���}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���}�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���}�j  sh�Kh�hRh�h�)��}�(h�}����}�j;  sh�K h�hRh�Nj0  h�)��}�(h�}����}�j>  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����}�j;  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�jh  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIje  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���}�je  sh�Kh�hRh�h�)��}�(h�}��P�}�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�}�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���}�h�)��}�(h�Kh�Kh�}����}�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����}�j�  sh�Kh�hRh�h�)��}�(h�}����}�j�  sh�K h�hRh�Nj0  h�)��}�(h�}����}�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����}�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�~�h�)��}�(h�Kh�Kh�}����~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�~�j�  sh�Kh�hRh�h�)��}�(h�}��P�~�j  sh�K h�hRh�Nj0  h�)��}�(h�}��P�~�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�~�j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�~�h�)��}�(h�Kh�Kh�}��P�~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�~�jI  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjF  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�~�jF  sh�Kh�hRh�h�)��}�(h�}����~�jg  sh�K h�hRh�Nj0  h�)��}�(h�}���~�jj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����~�jg  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���~�h�)��}�(h�Kh�Kh�}���~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����~�j�  sh�Kh�hRh�h�)��}�(h�}����~�j�  sh�K h�hRh�Nj0  h�)��}�(h�}����~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����~�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�~�h�)��}�(h�Kh�Kh�}���~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�~�j�  sh�Kh�hRh�h�)��}�(h�}����~�j�  sh�K h�hRh�Nj0  h�)��}�(h�}��P�~�j   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����~�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���~�h�)��}�(h�Kh�Kh�}���~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���~�j*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj'  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����~�j'  sh�Kh�hRh�h�)��}�(h�}����~�jH  sh�K h�hRh�Nj0  h�)��}�(h�}����~�jK  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����~�jH  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���~�h�)��}�(h�Kh�Kh�}��P�~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�~�ju  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjr  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����~�jr  sh�Kh�hRh�h�)��}�(h�}����~�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����~�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��~�h�)��}�(h�Kh�Kh�}����~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���~�j�  sh�Kh�hRh�h�)��}�(h�}���~�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���~�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���~�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���~�h�)��}�(h�Kh�Kh�}����~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����~�j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����~�j  sh�Kh�hRh�h�)��}�(h�}��P�~�j)  sh�K h�hRh�Nj0  h�)��}�(h�}��P�~�j,  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�~�j)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���~�h�)��}�(h�Kh�Kh�}���~�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���~�jV  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjS  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����~�jS  sh�Kh�hRh�h�)��}�(h�}����~�jt  sh�K h�hRh�Nj0  h�)��}�(h�}����~�jw  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����~�jt  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�� ��h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��� ��j�  sh�Kh�hRh�h�)��}�(h�}�����j�  sh�K h�hRh�Nj0  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�b�      j�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����j�  sh�Kh�hRh�h�)��}�(h�}��P��j
  sh�K h�hRh�Nj0  h�)��}�(h�}���
��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P��j
  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����j7  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj4  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����j4  sh�Kh�hRh�h�)��}�(h�}����jU  sh�K h�hRh�Nj0  h�)��}�(h�}��P��jX  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����jU  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��j  sh�Kh�hRh�h�)��}�(h�}��P��j�  sh�K h�hRh�Nj0  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��j�  sh�Kh�hRh�h�)��}�(h�}����j�  sh�K h�hRh�Nj0  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub� ��h�)��}�(h�Kh�Kh�}��&��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��&��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�� ��j  sh�Kh�hRh�h�)��}�(h�}���%��j6  sh�K h�hRh�Nj0  h�)��}�(h�}���$��j9  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���%��j6  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��'��h�)��}�(h�Kh�Kh�}���,��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���,��jc  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj`  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���'��j`  sh�Kh�hRh�h�)��}�(h�}��,��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���)��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��,��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�-��h�)��}�(h�Kh�Kh�}��3��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��3��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��-��j�  sh�Kh�hRh�h�)��}�(h�}���2��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���1��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���2��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��3��h�)��}�(h�Kh�Kh�}���9��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���9��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���3��j�  sh�Kh�hRh�h�)��}�(h�}��9��j  sh�K h�hRh�Nj0  h�)��}�(h�}��P5��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��9��j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}������h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}������jD  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjA  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������jA  sh�Kh�hRh�h�)��}�(h�}��;��jb  sh�K h�hRh�Nj0  h�)��}�(h�}��P>��je  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��;��jb  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P���h�)��}�(h�Kh�Kh�}���ǀ�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���ǀ�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P���j�  sh�Kh�hRh�h�)��}�(h�}��ǀ�j�  sh�K h�hRh�Nj0  h�)��}�(h�}��ƀ�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��ǀ�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PȀ�h�)��}�(h�Kh�Kh�}��P΀�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P΀�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PȀ�j�  sh�Kh�hRh�h�)��}�(h�}���̀�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���ɀ�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���̀�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�΀�h�)��}�(h�Kh�Kh�}��PԀ�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PԀ�j%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��΀�j"  sh�Kh�hRh�h�)��}�(h�}���Ӏ�jC  sh�K h�hRh�Nj0  h�)��}�(h�}��Ӏ�jF  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���Ӏ�jC  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��Հ�h�)��}�(h�Kh�Kh�}��ۀ�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��ۀ�jp  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjm  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���Հ�jm  sh�Kh�hRh�h�)��}�(h�}���ڀ�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���ـ�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���ڀ�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P܀�h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P܀�j�  sh�Kh�hRh�h�)��}�(h�}�����j�  sh�K h�hRh�Nj0  h�)��}�(h�}������j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��߀�h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���߀�j  sh�Kh�hRh�h�)��}�(h�}�����j$  sh�K h�hRh�Nj0  h�)��}�(h�}����j'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��jQ  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjN  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��jN  sh�Kh�hRh�h�)��}�(h�}�����jo  sh�K h�hRh�Nj0  h�)��}�(h�}�����jr  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����jo  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}��P���h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P���j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��j�  sh�Kh�hRh�h�)��}�(h�}�����j�  sh�K h�hRh�Nj0  h�)��}�(h�}�����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}������h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}������j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������j�  sh�Kh�hRh�h�)��}�(h�}�����j  sh�K h�hRh�Nj0  h�)��}�(h�}�����j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��A��h�)��}�(h�Kh�Kh�}���B��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���B��j2  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj/  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���A��j/  sh�Kh�hRh�h�)��}�(h�}��B��jP  sh�K h�hRh�Nj0  h�)��}�(h�}������jS  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��B��jP  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�D��h�)��}�(h�Kh�Kh�}��PI��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PI��j}  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjz  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��D��jz  sh�Kh�hRh�h�)��}�(h�}���H��j�  sh�K h�hRh�Nj0  h�)��}�(h�}��G��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���H��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��I��h�)��}�(h�Kh�Kh�}���O��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���O��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���I��j�  sh�Kh�hRh�h�)��}�(h�}��O��j�  sh�K h�hRh�Nj0  h�)��}�(h�}��PK��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��O��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}��V��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��V��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��j  sh�Kh�hRh�h�)��}�(h�}���U��j1  sh�K h�hRh�Nj0  h�)��}�(h�}���T��j4  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���U��j1  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��W��h�)��}�(h�Kh�Kh�}���\��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���\��j^  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj[  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���W��j[  sh�Kh�hRh�h�)��}�(h�}��P\��j|  sh�K h�hRh�Nj0  h�)��}�(h�}���[��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P\��j|  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��]��h�)��}�(h�Kh�Kh�}��Pc��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pc��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���]��j�  sh�Kh�hRh�h�)��}�(h�}���b��j�  sh�K h�hRh�Nj0  h�)��}�(h�}��^��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���b��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��c��h�)��}�(h�Kh�Kh�}��Pj��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pj��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���c��j�  sh�Kh�hRh�h�)��}�(h�}���i��j  sh�K h�hRh�Nj0  h�)��}�(h�}���h��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���i��j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��k��h�)��}�(h�Kh�Kh�}��p��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��p��j?  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj<  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���k��j<  sh�Kh�hRh�h�)��}�(h�}���o��j]  sh�K h�hRh�Nj0  h�)��}�(h�}���j��j`  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���o��j]  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��r��h�)��}�(h�Kh�Kh�}���v��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���v��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���r��j�  sh�Kh�hRh�h�)��}�(h�}��v��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���s��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��v��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Ps��h�)��}�(h�Kh�Kh�}���|��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���|��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Ps��j�  sh�Kh�hRh�h�)��}�(h�}��|��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���x��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��|��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��B��h�)��}�(h�Kh�Kh�}��PC��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PC��j   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���B��j  sh�Kh�hRh�h�)��}�(h�}���B��j>  sh�K h�hRh�Nj0  h�)��}�(h�}��A��jA  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���B��j>  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��D��h�)��}�(h�Kh�Kh�}��J��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��J��jk  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjh  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���D��jh  sh�Kh�hRh�h�)��}�(h�}���I��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���G��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���I��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�|�h�)��}�(h�Kh�Kh�}��\��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��\��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�|�j�  sh�Kh�hRh�h�)��}�(h�}���y�j�  sh�K h�hRh�Nj0  h�)��}�(h�}���dq�j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���y�j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�`��h�)��}�(h�Kh�Kh�}��b��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��b��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��`��j�  sh�Kh�hRh�h�)��}�(h�}���a��j  sh�K h�hRh�Nj0  h�)��}�(h�}���`��j"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���a��j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��`��h�)��}�(h�Kh�Kh�}��h��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��h��jL  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjI  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���`��jI  sh�Kh�hRh�h�)��}�(h�}���g��jj  sh�K h�hRh�Nj0  h�)��}�(h�}���f��jm  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���g��jj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��h��h�)��}�(h�Kh�Kh�}��Pn��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pn��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���h��j�  sh�Kh�hRh�h�)��}�(h�}���m��j�  sh�K h�hRh�Nj0  h�)��}�(h�}��j��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���m��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�r��h�)��}�(h�Kh�Kh�}��v��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��v��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��r��j�  sh�Kh�hRh�h�)��}�(h�}���u��j   sh�K h�hRh�Nj0  h�)��}�(h�}��p��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���u��j   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pw��h�)��}�(h�Kh�Kh�}��}��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��}��j-  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj*  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pw��j*  sh�Kh�hRh�h�)��}�(h�}���|��jK  sh�K h�hRh�Nj0  h�)��}�(h�}���w��jN  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���|��jK  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�C��h�)��}�(h�Kh�Kh�}���C��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���C��jx  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIju  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��C��ju  sh�Kh�hRh�h�)��}�(h�}��PC��j�  sh�K h�hRh�Nj0  h�)��}�(h�}����j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PC��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�D��h�)��}�(h�Kh�Kh�}���I��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���I��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��D��j�  sh�Kh�hRh�h�)��}�(h�}��PI��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���E��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PI��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�K��h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��K��j  sh�Kh�hRh�h�)��}�(h�}���O��j,  sh�K h�hRh�Nj0  h�)��}�(h�}���L��j/  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���O��j,  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��R��h�)��}�(h�Kh�Kh�}��PV��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PV��jY  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjV  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���R��jV  sh�Kh�hRh�h�)��}�(h�}���U��jw  sh�K h�hRh�Nj0  h�)��}�(h�}���S��jz  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���U��jw  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�S��h�)��}�(h�Kh�Kh�}���\��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���\��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��S��j�  sh�Kh�hRh�h�)��}�(h�}��\��j�  sh�K h�hRh�Nj0  h�)��}�(h�}���Y��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��\��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�_��h�)��}�(h�Kh�Kh�}���b��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���b��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��_��j�  sh�Kh�hRh�h�)��}�(h�}��Pb��j  sh�K h�hRh�Nj0  h�)��}�(h�}��`��j  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Pb��j  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pd��h�)��}�(h�Kh�Kh�}��Pi��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pi��j:  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj7  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pd��j7  sh�Kh�hRh�h�)��}�(h�}���h��jX  sh�K h�hRh�Nj0  h�)��}�(h�}���f��j[  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���h��jX  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��k��h�)��}�(h�Kh�Kh�}��p��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��p��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���k��j�  sh�Kh�hRh�h�)��}�(h�}���o��j�  sh�K h�hRh�Nj0  h�)��}�(h�}��k��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���o��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��o��h�)��}�(h�Kh�Kh�}��Pv��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pv��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���o��j�  sh�Kh�hRh�h�)��}�(h�}���u��j�  sh�K h�hRh�Nj0  h�)��}�(h�}��u��j�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���u��j�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��x��h�)��}�(h�Kh�Kh�}��}��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��}��j   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���x��j   sh�Kh�hRh�h�)��}�(h�}���|��j9   sh�K h�hRh�Nj0  h�)��}�(h�}���z��j<   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���|��j9   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��B��h�)��}�(h�Kh�Kh�}��PC��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PC��jf   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjc   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���B��jc   sh�Kh�hRh�h�)��}�(h�}���B��j�   sh�K h�hRh�Nj0  h�)��}�(h�}���~��j�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���B��j�   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�D��h�)��}�(h�Kh�Kh�}���I��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���I��j�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��D��j�   sh�Kh�hRh�h�)��}�(h�}��PI��j�   sh�K h�hRh�Nj0  h�)��}�(h�}��PE��j�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PI��j�   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PL��h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��j�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PL��j�   sh�Kh�hRh�h�)��}�(h�}���O��j!  sh�K h�hRh�Nj0  h�)��}�(h�}��PM��j!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���O��j!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PU��h�)��}�(h�Kh�Kh�}��PV��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PV��jG!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjD!  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PU��jD!  sh�Kh�hRh�h�)��}�(h�}���U��je!  sh�K h�hRh�Nj0  h�)��}�(h�}��R��jh!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���U��je!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��V��h�)��}�(h�Kh�Kh�}���\��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���\��j�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�!  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���V��j�!  sh�Kh�hRh�h�)��}�(h�}��\��j�!  sh�K h�hRh�Nj0  h�)��}�(h�}��PX��j�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��\��j�!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�]��h�)��}�(h�Kh�Kh�}��c��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��c��j�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�!  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��]��j�!  sh�Kh�hRh�h�)��}�(h�}���b��j�!  sh�K h�hRh�Nj0  h�)��}�(h�}���a��j�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���b��j�!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�d��h�)��}�(h�Kh�Kh�}���i��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���i��j("  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj%"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��d��j%"  sh�Kh�hRh�h�)��}�(h�}��i��jF"  sh�K h�hRh�Nj0  h�)��}�(h�}��Pe��jI"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��i��jF"  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��i��h�)��}�(h�Kh�Kh�}���o��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���o��js"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjp"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���i��jp"  sh�Kh�hRh�h�)��}�(h�}��o��j�"  sh�K h�hRh�Nj0  h�)��}�(h�}��Pn��j�"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��o��j�"  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pp��h�)��}�(h�Kh�Kh�}��v��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��v��j�"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pp��j�"  sh�Kh�hRh�h�)��}�(h�}���u��j�"  sh�K h�hRh�Nj0  h�)��}�(h�}���q��j�"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���u��j�"  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��v��h�)��}�(h�Kh�Kh�}���|��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���|��j	#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���v��j#  sh�Kh�hRh�h�)��}�(h�}��|��j'#  sh�K h�hRh�Nj0  h�)��}�(h�}��Pw��j*#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��|��j'#  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��B��h�)��}�(h�Kh�Kh�}��D��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��D��jT#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjQ#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���B��jQ#  sh�Kh�hRh�h�)��}�(h�}���C��jr#  sh�K h�hRh�Nj0  h�)��}�(h�}���}��ju#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���C��jr#  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PA��h�)��}�(h�Kh�Kh�}��PJ��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PJ��j�#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PA��j�#  sh�Kh�hRh�h�)��}�(h�}���I��j�#  sh�K h�hRh�Nj0  h�)��}�(h�}��PE��j�#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���I��j�#  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��K��h�)��}�(h�Kh�Kh�}��PQ��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PQ��j�#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���K��j�#  sh�Kh�hRh�h�)��}�(h�}���P��j$  sh�K h�hRh�Nj0  h�)��}�(h�}���O��j$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���P��j$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��S��h�)��}�(h�Kh�Kh�}��PW��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PW��j5$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj2$  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���S��j2$  sh�Kh�hRh�h�)��}�(h�}���V��jS$  sh�K h�hRh�Nj0  h�)��}�(h�}���T��jV$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���V��jS$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��S��h�)��}�(h�Kh�Kh�}���]��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���]��j�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj}$  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���S��j}$  sh�Kh�hRh�h�)��}�(h�}��]��j�$  sh�K h�hRh�Nj0  h�)��}�(h�}��P\��j�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��]��j�$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�^��h�)��}�(h�Kh�Kh�}���c��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���c��j�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�$  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��^��j�$  sh�Kh�hRh�h�)��}�(h�}��Pc��j�$  sh�K h�hRh�Nj0  h�)��}�(h�}���_��j�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Pc��j�$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�e��h�)��}�(h�Kh�Kh�}��Pj��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pj��j%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��e��j%  sh�Kh�hRh�h�)��}�(h�}���i��j4%  sh�K h�hRh�Nj0  h�)��}�(h�}��i��j7%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���i��j4%  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�l��h�)��}�(h�Kh�Kh�}��Pq��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pq��ja%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj^%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��l��j^%  sh�Kh�hRh�h�)��}�(h�}���p��j%  sh�K h�hRh�Nj0  h�)��}�(h�}��o��j�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���p��j%  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��r��h�)��}�(h�Kh�Kh�}���w��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���w��j�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���r��j�%  sh�Kh�hRh�h�)��}�(h�}��Pw��j�%  sh�K h�hRh�Nj0  h�)��}�(h�}���v��j�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Pw��j�%  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��z��h�)��}�(h�Kh�Kh�}��P~��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P~��j�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���z��j�%  sh�Kh�hRh�h�)��}�(h�}���}��j&  sh�K h�hRh�Nj0  h�)��}�(h�}��Pz��j&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���}��j&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}��PŇ�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PŇ�jB&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj?&  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������j?&  sh�Kh�hRh�h�)��}�(h�}���ć�j`&  sh�K h�hRh�Nj0  h�)��}�(h�}��ć�jc&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���ć�j`&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Ƈ�h�)��}�(h�Kh�Kh�}���ˇ�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���ˇ�j�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�&  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Ƈ�j�&  sh�Kh�hRh�h�)��}�(h�}��ˇ�j�&  sh�K h�hRh�Nj0  h�)��}�(h�}���Ƈ�j�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��ˇ�j�&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��̇�h�)��}�(h�Kh�Kh�}��P҇�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P҇�j�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�&  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubs�       h�Kh�hRh�h�)��}�(h�Kh�Kh�}���̇�j�&  sh�Kh�hRh�h�)��}�(h�}���ч�j�&  sh�K h�hRh�Nj0  h�)��}�(h�}��·�j�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���ч�j�&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��Ӈ�h�)��}�(h�Kh�Kh�}��ه�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��ه�j#'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj '  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���Ӈ�j '  sh�Kh�hRh�h�)��}�(h�}���؇�jA'  sh�K h�hRh�Nj0  h�)��}�(h�}���ׇ�jD'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���؇�jA'  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PՇ�h�)��}�(h�Kh�Kh�}���߇�h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���߇�jn'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjk'  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PՇ�jk'  sh�Kh�hRh�h�)��}�(h�}��P߇�j�'  sh�K h�hRh�Nj0  h�)��}�(h�}��Pۇ�j�'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P߇�j�'  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����j�'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�'  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������j�'  sh�Kh�hRh�h�)��}�(h�}�����j�'  sh�K h�hRh�Nj0  h�)��}�(h�}�����j�'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j�'  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}��P��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��j(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��j(  sh�Kh�hRh�h�)��}�(h�}�����j"(  sh�K h�hRh�Nj0  h�)��}�(h�}�����j%(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����j"(  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����jO(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjL(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����jL(  sh�Kh�hRh�h�)��}�(h�}��P��jm(  sh�K h�hRh�Nj0  h�)��}�(h�}�����jp(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P��jm(  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��h�)��}�(h�Kh�Kh�}��P���h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P���j�(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��j�(  sh�Kh�hRh�h�)��}�(h�}������j�(  sh�K h�hRh�Nj0  h�)��}�(h�}�����j�(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}������j�(  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}������h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}������j�(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������j�(  sh�Kh�hRh�h�)��}�(h�}��P���j)  sh�K h�hRh�Nj0  h�)��}�(h�}������j)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P���j)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����h�)��}�(h�Kh�Kh�}������h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}������j0)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj-)  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����j-)  sh�Kh�hRh�h�)��}�(h�}������jN)  sh�K h�hRh�Nj0  h�)��}�(h�}��Ё��jQ)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}������jN)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����j{)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjx)  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������jx)  sh�Kh�hRh�h�)��}�(h�}������j�)  sh�K h�hRh�Nj0  h�)��}�(h�}��Ј��j�)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}������j�)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���_�h�)��}�(h�Kh�Kh�}��Ў��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Ў��j�)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�)  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����_�j�)  sh�Kh�hRh�h�)��}�(h�}��Г��j�)  sh�K h�hRh�Nj0  h�)��}�(h�}��В��j�)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Г��j�)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����j*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj*  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����j*  sh�Kh�hRh�h�)��}�(h�}������j/*  sh�K h�hRh�Nj0  h�)��}�(h�}������j2*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}������j/*  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����h�)��}�(h�Kh�Kh�}��А��h�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��А��j\*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjY*  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������jY*  sh�Kh�hRh�h�)��}�(h�}��P���jz*  sh�K h�hRh�Nj0  h�)��}�(h�}�����j}*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P���jz*  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ubuh�Kh�hRh�Nj0  h�h�hhK ��h��R�(KKK��h!�CH      Y@        �8��8V�@             xz@9��8��I@                      �?�t�bubsh�Kh�hRj�  h�hIh�j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�K h�hRj�  hhK ��h��R�(KKK��h!�C �������?(\���(�?�������?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bub�_originalPosition�h�)��}�(h�}�h�Kh�hRj�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bub�_aspect�h7�_adjustable��box��_anchor��C��_stale_viewlims�}�(h~�h��u�_sharex�N�_sharey�h>�bbox�h��dataLim�h�)��}�(h�}�h�Kh�hRj�  hhK ��h��R�(KKK��h!�C         ���`C!�     �E@ڜ��H��?�t�bj�  hhK ��h��R�(KK��h!�C      �?�>���q?�t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �      �      ��      ���t�bub�_viewLim�j	  �
transScale�j�  �	transAxes�h��transLimits�j	  �	transData�h��_xaxis_transform�h��_yaxis_transform�j	  �_subplotspec�N�_box_aspect�N�_axes_locator��$mpl_toolkits.axes_grid1.axes_divider��AxesLocator���)��}�(�_axes_divider�j+  �AxesDivider���)��}�(hBh>�_xref��!mpl_toolkits.axes_grid1.axes_size��AxesX���)��}�(hBh>j�*  G?�      �_ref_ax�Nub�_yref�j+  �AxesY���)��}�(hBh>j�*  G?�      j+  Nub�_fig�hG�_pos�N�_horizontal�]�(j+  j+  �Fixed���)��}��
fixed_size�G?�������sbj+  )��}�j +  Ksbe�	_vertical�]�j+  aj�*  j�*  j�*  N�
_xrefindex�K �
_yrefindex�K �_locator�Nub�_nx�K�_ny�K �_nx1�K�_ny1�Kub�	_children�]�(�matplotlib.patches��	Rectangle���)��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQ�
_nolegend_�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx��_hatch_color�(G        G        G        G?�      t��_fill���_original_edgecolor�N�
_edgecolor�(G        G        G        G        t��_original_facecolor�hhK ��h��R�(KK��h!�C �?�������?TTTTTT�?      �?�t�b�
_facecolor�(G?�G?ܜ�����G?�TTTTTTG?�      t��
_linewidth�G?�333333�_unscaled_dash_pattern�K N���_dash_pattern�G        N���
_linestyle��solid��_antialiased���_hatch�N�	_capstyle��matplotlib._enums��CapStyle����butt���R��
_joinstyle�j\+  �	JoinStyle����miter���R��_x0�j?+  �_y0�h0h!C���`C!⿔��R��_width�h0h!C       @���R��_height�h0h!C@����[�?���R��angle�G        �_rotation_point��xy��_aspect_ratio_correction�G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj[  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�+  ji+  h0h!Cr��id^῔��R�jm+  h0h!C        ���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�+  ji+  h0h!C�iLr��࿔��R�jm+  h0h!C      �?���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�+  ji+  h0h!C�H0�L�߿���R�jm+  h0h!C        ���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj<  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�+  ji+  h0h!C	���+޿���R�jm+  h0h!C      �?���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�+  ji+  h0h!C3_ѥܿ���R�jm+  h0h!C       @���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j,  ji+  h0h!C$��* ۿ���R�jm+  h0h!C      @���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j4,  ji+  h0h!C0�<U�ٿ���R�jm+  h0h!C      @���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjh  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jQ,  ji+  h0h!C;�%N�ؿ���R�jm+  h0h!C      @���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jn,  ji+  h0h!CI�_ֿَ���R�jm+  h0h!C        ���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�,  ji+  h0h!CV|Tq	տ���R�jm+  h0h!C       @���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjI  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�,  ji+  h0h!Ca��]�ӿ���R�jm+  h0h!C      @���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�,  ji+  h0h!Cof����ѿ���R�jm+  h0h!C      @���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�,  ji+  h0h!Cz���wп���R�jm+  h0h!C      *@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj*  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�,  ji+  h0h!C�doG�Ϳ���R�jm+  h0h!C      &@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNju  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j-  ji+  h0h!C'�����ʿ���R�jm+  h0h!C       @���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j9-  ji+  h0h!CAuµO�ǿ���R�jm+  h0h!C      &@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jV-  ji+  h0h!C\_����Ŀ���R�jm+  h0h!C      3@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjV  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  js-  ji+  h0h!CsI �W������R�jm+  h0h!C      4@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�-  ji+  h0h!Cg�>�U�����R�jm+  h0h!C      >@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�-  ji+  h0h!CJ;���>�����R�jm+  h0h!C      :@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj7  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�-  ji+  h0h!C�Z��'�����R�jm+  h0h!C      ?@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�-  ji+  h0h!C`�o#�!�����R�jm+  h0h!C      E@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j.  ji+  h0h!C��V`e瓿���R�jm+  h0h!C     �E@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j!.  ji+  h0h!C�>���q?���R�jm+  h0h!C      >@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjc  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j>.  ji+  h0h!C�~�lXМ?���R�jm+  h0h!C      <@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j[.  ji+  h0h!C�����?���R�jm+  h0h!C      4@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jx.  ji+  h0h!CP�r�b�?���R�jm+  h0h!C      6@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjD  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�.  ji+  h0h!C #H�x�?���R�jm+  h0h!C      =@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�.  ji+  h0h!C�N����?���R�jm+  h0h!C      5@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�.  ji+  h0h!C`��]v��?���R�jm+  h0h!C      2@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj%  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�.  ji+  h0h!CD�}:���?���R�jm+  h0h!C      1@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjp  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j	/  ji+  h0h!C,�Nn��?���R�jm+  h0h!C      ,@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j&/  ji+  h0h!C�����?���R�jm+  h0h!C      (@���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jC/  ji+  h0h!C���e�?���R�jm+  h0h!C      *@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjQ  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j`/  ji+  h0h!Cp��p�?���R�jm+  h0h!C        ���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j}/  ji+  h0h!Cd�I�.��?���R�jm+  h0h!C      &@���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�/  ji+  h0h!CX+����?���R�jm+  h0h!C      �?���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj2  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�/  ji+  h0h!CJ�����?���R�jm+  h0h!C      @���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj}  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�/  ji+  h0h!C>A��h�?���R�jm+  h0h!C      �?���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�/  ji+  h0h!C2��~&��?���R�jm+  h0h!C       @���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j0  ji+  h0h!C$WTm�(�?���R�jm+  h0h!C      �?���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj^  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j+0  ji+  h0h!C�[���?���R�jm+  h0h!C       @���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jH0  ji+  h0h!Cm%J`4�?���R�jm+  h0h!C      �?���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  je0  ji+  h0h!C ��8��?���R�jm+  h0h!C        ���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj?  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�0  ji+  h0h!CzA{��?���R�jm+  h0h!C        ���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�0  ji+  h0h!C�
���?���R�jm+  h0h!C      �?���R�jq+  h0h!C ����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�0  ji+  h0h!Cl�����?���R�jm+  h0h!C        ���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj   hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�0  ji+  h0h!C���h�?���R�jm+  h0h!C      �?���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjk  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  jL+  jP+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�0  ji+  h0h!C`WL�i+�?���R�jm+  h0h!C      �?���R�jq+  h0h!C@����[�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  hhK ��h��R�(KK��h!�C �������?xxxxxx�?�������?      �?�t�bjP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j1  ji+  h0h!C(�R�J߿���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j61  ji+  h0h!COajJ��ݿ���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjL  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jS1  ji+  h0h!Ctځ���ܿ���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jp1  ji+  h0h!C�S�A]ۿ���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�1  ji+  h0h!C�̰|�%ڿ���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj-  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�1  ji+  h0h!C�E���ؿ���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjx  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�1  ji+  h0h!C��H7�׿���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�1  ji+  h0h!C68���ֿ���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j2  ji+  h0h!C\��Hտ���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjY  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j2  ji+  h0h!C�*&{-Կ���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j;2  ji+  h0h!C��=���ҿ���R�jm+  h0h!C       @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jX2  ji+  h0h!C�UG|�ѿ���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj:  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  ju2  ji+  h0h!C��l�#kп���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�2  ji+  h0h!C<'�gο���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�2  ji+  h0h!C�7���˿���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj   hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�2  ji+  h0h!C�f�3�ɿ���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjf   hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�2  ji+  h0h!C"����ǿ���R�jm+  h0h!C       @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�   hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j3  ji+  h0h!Cp��WѬĿ���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�   hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j#3  ji+  h0h!C���# >¿���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjG!  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j@3  ji+  h0h!C�C�ݞ�����R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�!  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j]3  ji+  h0h!C�|�x{������R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�!  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jz3  ji+  h0h!CHa�䵿���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj("  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�3  ji+  h0h!C�E]�������R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjs"  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�3  ji+  h0h!C�Tv��R�����R�jm+  h0h!C       @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�"  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�3  ji+  h0h!C`<dh�/�����R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj	#  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�3  ji+  h0h!C����{t�����R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjT#  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j4  ji+  h0h!C�=Y��v�?���R�jm+  h0h!C      $@���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�#  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j(4  ji+  h0h!C`5s�0�?���R�jm+  h0h!C       @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�#  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jE4  ji+  h0h!C �ވ/S�?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj5$  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jb4  ji+  h0h!C�y,��?���R�jm+  h0h!C       @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�$  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j4  ji+  h0h!CP���\�?���R�jm+  h0h!C       @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�$  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�4  ji+  h0h!C��U����?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj%  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�4  ji+  h0h!C��b!��?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNja%  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�4  ji+  h0h!C��L�A>�?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�%  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�4  ji+  h0h!Cp��?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�%  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j5  ji+  h0h!C$�L��?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjB&  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j-5  ji+  h0h!C���U��?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�&  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jJ5  ji+  h0h!C�*����?���R�jm+  h0h!C      @���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�&  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jg5  ji+  h0h!C<8b�g�?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj#'  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�5  ji+  h0h!C���4k�?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjn'  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�5  ji+  h0h!C�)(���?���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�'  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�5  ji+  h0h!C�������?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj(  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�5  ji+  h0h!C�7�[>�?���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjO(  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�5  ji+  h0h!C^����H�?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�(  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j6  ji+  h0h!C8E����?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�(  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j26  ji+  h0h!C̌)H��?���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj0)  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jO6  ji+  h0h!C�Ruà��?���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj{)  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  jl6  ji+  h0h!C��]]�%�?���R�jm+  h0h!C        ���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�)  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�6  ji+  h0h!C�`F�Q]�?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj*  hONhP�hQj3+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jC+  jD+  jE+  �jF+  NjG+  jH+  jI+  j1  jP+  (G?�������G?�xxxxxxG?�������G?�      t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  j�6  ji+  h0h!Cv�.����?���R�jm+  h0h!C      �?���R�jq+  h0h!C�m���u�?���R�ju+  G        jv+  jw+  jx+  G?�      ub�matplotlib.lines��Line2D���)��}�(h@�hANhBh�hChGhIj	  hJ�hK�hL�hMNhNj\*  hONhP�hQ�	_child100�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j-+  �remove���R�hjNhkNhlNhmNhnhohphs]�]�����hx��_dashcapstyle�ja+  �_dashjoinstyle�jd+  �round���R��_solidjoinstyle�j�6  �_solidcapstyle�j^+  j�6  ��R��_linestyles�N�
_drawstyle��default�jR+  G?�      jS+  K N��jU+  G        N��jW+  �-��	_invalidx���_color��#111111��_marker��matplotlib.markers��MarkerStyle���)��}�(�_marker_function�h�j�6  �_set_nothing���R��_user_transform�N�_user_capstyle�N�_user_joinstyle�N�
_fillstyle��full�j�6  �None�j#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�C �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nub�	_alt_path�N�_alt_transform�N�_snap_threshold�Njb+  j�6  j[+  ja+  �_filled��ub�	_gapcolor�N�
_markevery�N�_markersize�G@      jY+  ��_markeredgecolor��auto��_markeredgewidth�G        �_markerfacecolor��auto��_markerfacecoloralt��none��	_invalidy���_pickradius�K�
ind_offset�K �_xorig�]�(K Ke�_yorig�]�(K K ej�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�b�_xy�hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  j>  j5  j;  �	_subslice���	_x_filled�Nube�
_colorbars�]��spines��matplotlib.spines��Spines���)��}�(�left�j"7  �Spine���)��}�(h@�hANhBh�hChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  (G?陙����G?陙����G?陙����G?�      t�jE+  �jF+  �.8�jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j^+  �
projecting���R�jb+  jg+  �
spine_type�j'7  �axis��matplotlib.axis��YAxis���)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj?  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx��_remove_overlapping_locs���isDefault_label���major�j>7  �Ticker���)��}�(j'+  �matplotlib.ticker��AutoLocator���)��}�(�_nbins�h7�
_symmetric���_prune�N�_min_n_ticks�K�_steps�hhK ��h��R�(KK��h!�C(      �?       @      @      @      $@�t�b�_extended_steps�hhK ��h��R�(KK
��h!�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�b�_integer��j=7  j@7  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jL7  �jM7  �jN7  jQ7  �minor�jP7  )��}�(j'+  jS7  �NullLocator���)��}�j=7  jk7  sb�
_formatter�jS7  �NullFormatter���)��}�(j=7  jk7  �locs�hhK ��h��R�(KK ��h!�j�6  t�bub�_locator_is_default���_formatter_is_default��ubhchZ)��}�(h]]��units�ah`hbhc}�j�7  }�K �	functools��partial���h�h>�_unit_change_handler���R���R�(j�7  h���}��event��builtins��object���)��sNt�bssheKhfNhg��(K �ub�_autolabelpos���label��matplotlib.text��Text���)��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  h0h!C������7@���R�j�  G?�      �_text��	Residuals�j�6  �.15��_fontproperties��matplotlib.font_manager��FontProperties���)��}�(�_family�]��
sans-serif�a�_slant��normal��_variant��normal��_weight��normal��_stretch��normal��_file�N�_size�G@&      �_math_fontfamily��
dejavusans�ub�_usetex���_parse_math���_wrap���_verticalalignment��bottom��_horizontalalignment��center��_multialignment�N�	_rotation�G@V�     �_transform_rotates_text���_bbox_patch�N�	_renderer�N�_linespacing�G?�333333�_rotation_mode��anchor�ub�
offsetText�j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  h0h!Cr�q�}@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  �      j�7  j�7  j�7  j�7  �normal�j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  �baseline�j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nub�labelpad�G@      j7  K�_major_tick_kw�}�(�gridOn���tick1On���tick2On���label1On���label2On��u�_minor_tick_kw�}�(j�7  �j�7  �j�7  �j�7  �j�7  �u�label_position�j'7  �offset_text_position�j'7  �_scale��matplotlib.scale��LinearScale���)���	converter�Nj�7  N�_autoscale_on���zorder�G?�      �
majorTicks�]�(j>7  �YTick���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj#  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx��_loc�h0h!C������鿔��R��_major��j�7  G        jm+  G?�      �	_base_pad�G@      �_labelrotation�j�6  K ���_zorder�G@ z�G��	tick1line�j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  �None�j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j)8  �_set_tickleft���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j8  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nub�	tick2line�j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jO8  �_set_tickright���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j8  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nub�gridline�j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�jm8  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j8  ��j7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nub�label1�j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j8  j�7  �−0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  �center_baseline�j�7  �right�j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nub�label2�j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j8  j�7  j�8  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nub�_tickdir��out��_pad�G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333㿔��R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�8  j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�8  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C433333㿔t�bj7  hhK ��h��R�(KKK��h!�C        433333㿔t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        433333㿔t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j 9  jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�8  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j9  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�8  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�433333㿔t�bj7  hhK ��h��R�(KKK��h!�C         433333�      �?433333㿔t�bj#  j�  j5  j�  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�8  j�7  �−0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�8  j�7  jB9  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ٿ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j_9  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C        ������ٿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        ������ٿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j_9  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j_9  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ٿ������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ٿ      �?������ٿ�t�bj#  j
  j5  j  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j_9  j�7  �−0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j_9  j�7  j�9  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ɿ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j:  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C        ������ɿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        ������ɿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j:  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j:  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ɿ������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ɿ      �?������ɿ�t�bj#  j  j5  j  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j:  j�7  �−0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j:  j�7  j�:  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C        ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�:  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C                �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�:  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�:  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�bj7  hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  j(  j5  j%  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�:  j�7  �0.0�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�:  j�7  jj;  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�;  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C        �������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�;  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�;  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  j7  j5  j4  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�;  j�7  �0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�;  j�7  j"<  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j?<  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C        �������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j?<  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j?<  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  jF  j5  jC  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j?<  j�7  �0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j?<  j�7  j�<  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333�?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�<  ��j7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C433333�?�t�bj7  hhK ��h��R�(KKK��h!�C        433333�?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        433333�?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�<  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�<  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�?433333�?�t�bj7  hhK ��h��R�(KKK��h!�C         433333�?      �?433333�?�t�bj#  jU  j5  jR  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�<  j�7  �0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�<  j�7  j�=  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j&8  jU+  j'8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�=  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jM8  jU+  jN8  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�=  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jk8  jU+  jl8  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�=  ��j7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�=  j�7  �0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�=  j�7  j4>  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ube�
minorTicks�]�j8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj7  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        jm+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j_>  j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�K aj7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j{>  jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�Kaj7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjv  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�>  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  ]�(K K ej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@333333ubaububj}7  jS7  �ScalarFormatter���)��}�(�_offset_threshold�K�offset�K �
_useOffset��j�7  ��_useMathText���orderOfMagnitude�K �format��%1.1f��_scientific���_powerlimits�]�(J����Ke�
_useLocale��j=7  jk7  j�7  hhK ��h��R�(KK	��h!�CH�������433333㿚�����ٿ������ɿ        �������?�������?433333�?�������?�t�bubj�7  �j�7  �ubjv7  jw7  hchZ)��}�(h]]�j�7  ah`hbhc}�j�7  }�K j�7  h�h�j�7  ��R���R�(j�>  h���}�j�7  j�7  )��sNt�bssheKhfNhg��(K �ubj�7  �j�7  j�7  )��}�(h@�hANhBNhChGhIjS	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  h0h!C�q�)�@���R�j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@&      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G@V�     j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�7  ubj�7  j�7  )��}�(h@�hANhBNhChGhIj_	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  h0h!Cr�q�}@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�7  G@      j7  Kj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  j'7  j�7  j'7  j�7  j�7  j�7  Nj�7  Nj 8  �j8  G?�      j8  ]�(j8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj~  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������鿔��R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j2?  j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j#?  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jN?  jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j#?  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�jj?  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j#?  ��j7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j#?  j�7  �−0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j#?  j�7  j�?  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333㿔��R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�?  j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�?  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�?  jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�?  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C433333㿔t�bj7  hhK ��h��R�(KKK��h!�C      �?433333㿔t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?433333㿔t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNjG  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j@  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�?  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�433333㿔t�bj7  hhK ��h��R�(KKK��h!�C         433333�      �?433333㿔t�bj#  jM  j5  jJ  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�?  j�7  �−0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�?  j�7  j8@  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ٿ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  jU@  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  jU@  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C      �?������ٿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?������ٿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  jU@  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ٿ������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ٿ      �?������ٿ�t�bj#  j\  j5  jY  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  jU@  j�7  �−0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  jU@  j�7  j�@  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ɿ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  jA  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  jA  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C      �?������ɿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?������ɿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  jA  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ɿ������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ɿ      �?������ɿ�t�bj#  jk  j5  jh  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  jA  j�7  �−0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  jA  j�7  j�A  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C        ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�A  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�A  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�A  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�bj7  hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  jz  j5  jw  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�A  j�7  �0.0�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�A  j�7  j`B  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j}B  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j}B  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j}B  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  j�  j5  j�  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j}B  j�7  �0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j}B  j�7  jC  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j5C  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j5C  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j5C  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  j�  j5  j�  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j5C  j�7  �0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j5C  j�7  j�C  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333�?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�C  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�C  ��j7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C433333�?�t�bj7  hhK ��h��R�(KKK��h!�C      �?433333�?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?433333�?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj_8  j�6  �      )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�C  ��j7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�?433333�?�t�bj7  hhK ��h��R�(KKK��h!�C         433333�?      �?433333�?�t�bj#  j�  j5  j�  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�C  j�7  �0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�C  j�7  j�D  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j0?  jU+  j1?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�K aj7  j�D  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jL?  jU+  jM?  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  ]�Kaj7  j�D  ��j7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jh?  jU+  ji?  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  j�D  ��j7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�D  j�7  �0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�D  j�7  j*E  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubejD>  ]�j8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        jm+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jTE  j+8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�K aj7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jpE  jQ8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j.8  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�Kaj7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�E  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K Kej7  ]�(K K ej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj-  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj4  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@333333ubaubj8  G@      �_bounds�Nh��outward�G        ��j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C         ����p�        �J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ub�_patch_type��line��_patch_transform�j�  )��}�(h�}�h�Kh�hRh�Nububj�8  j)7  )��}�(h@�hANhBh�hChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  j�8  j=7  jA7  j8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?����p�      �?�J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububj�7  j)7  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  j�7  j=7  j>7  �XAxis���)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�	  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jL7  �jM7  �jN7  jP7  )��}�(j'+  jU7  )��}�(jX7  h7jY7  �jZ7  Nj[7  Kj\7  hhK ��h��R�(KK��h!�C(      �?       @      @      @      $@�t�bjc7  hhK ��h��R�(KK
��h!�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�bjj7  �j=7  j�E  ubj}7  j�>  )��}�(j�>  Kj�>  K j�>  �j�7  �j�>  �j�>  K j�>  �%1.0f�j�>  �j�>  j�>  j�>  �j=7  j�E  j�7  hhK ��h��R�(KK��h!�C              9@      I@�t�bubj�7  �j�7  �ubjv7  jP7  )��}�(j'+  jz7  )��}�j=7  j�E  sbj}7  j7  )��}�(j=7  j�E  j�7  hhK ��h��R�(KK ��h!�j�6  t�bubj�7  �j�7  �ubhchZ)��}�(h]]�j�7  ah`hbhc}�j�7  }�K j�7  h�h�j�7  ��R���R�(j2F  h~��}�j�7  j�7  )��sNt�bssheKhfNhg��(K �ubj�7  �j�7  j�7  )��}�(h@�hANhBNhChGhIjk	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  h0h!C      8@���R�j�7  �Distribution�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@&      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  �top�j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�7  j�7  )��}�(h@�hANhBNhChGhIjw	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  h0h!C9��8�c9@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�7  G@      j7  Kj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  j�7  j�7  j�7  j�7  j�7  )��j�7  Nj�7  Nj 8  �j8  G?�      j8  ]�(j>7  �XTick���)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�	  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C        ���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j~F  �_set_tickdown���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  joF  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C                �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�F  �_set_tickup���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  joF  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�F  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  joF  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  joF  j�  K j�7  �0�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  joF  j�  Kj�7  jG  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNjC
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      9@���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j0G  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j!G  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      9@�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      9@        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      9@        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jfG  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j!G  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�G  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j!G  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j!G  j�  K j�7  �25�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j!G  j�  Kj�7  j�G  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      I@���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j|F  jU+  j}F  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�G  ��j7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�F  jU+  j�F  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�G  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�F  jU+  j�F  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j�G  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�G  j�  K j�7  �50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�G  j�  Kj�7  jNH  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubejD>  ]�jaF  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        jm+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jxH  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�K aj7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�H  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�K aj7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj   hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�H  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K K ej7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  Kj�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@333333uba�_tick_position�j�7  ubj8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                 33333�F@        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�NububjKF  j)7  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  jKF  j=7  j�E  j8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?33333�F@      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububub�xaxis�j�E  �yaxis�jA7  jP+  �white��_frameon���
_axisbelow���_rasterization_zorder�N�ignore_existing_data_limits��hchZ)��}�(h]]�(�xlim_changed��ylim_changed��zlim_changed�eh`hbhc}�heK hfNhg��ub�_xmargin�G?��������_ymargin�G?��������_tight�N�_use_sticky_edges���
_get_lines��matplotlib.axes._base��_process_plot_var_args���)��}�(�axes�h��command��plot�ub�_get_patches_for_fill�j#I  )��}�(j&I  h�j'I  �fill�ub�_gridOn���_mouseover_set�hX�_OrderedSet���)��}��_od��collections��OrderedDict���)R�sb�
child_axes�]��_current_image�N�_projection_init�N�legend_�N�
containers�]�(�matplotlib.container��BarContainer���(j1+  jy+  j�+  j�+  j�+  j�+  j
,  j',  jD,  ja,  j~,  j�,  j�,  j�,  j�,  j-  j,-  jI-  jf-  j�-  j�-  j�-  j�-  j�-  j.  j1.  jN.  jk.  j�.  j�.  j�.  j�.  j�.  j/  j6/  jS/  jp/  j�/  j�/  j�/  j�/  j0  j0  j;0  jX0  ju0  j�0  j�0  j�0  j�0  t�����}�(�patches�]�(j1+  jy+  j�+  j�+  j�+  j�+  j
,  j',  jD,  ja,  j~,  j�,  j�,  j�,  j�,  j-  j,-  jI-  jf-  j�-  j�-  j�-  j�-  j�-  j.  j1.  jN.  jk.  j�.  j�.  j�.  j�.  j�.  j/  j6/  jS/  jp/  j�/  j�/  j�/  j�/  j0  j0  j;0  jX0  ju0  j�0  j�0  j�0  j�0  e�errorbar�N�
datavalues�hhK ��h��R�(KK2��h!�B�         @              �?              �?       @      @      @      @               @      @      @      *@      &@       @      &@      3@      4@      >@      :@      ?@      E@     �E@      >@      <@      4@      6@      =@      5@      2@      1@      ,@      (@      *@              &@      �?      @      �?       @      �?       @      �?                      �?              �?      �?�t�b�orientation��
horizontal�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j>I  �remove���R�hQ�_container0��stale��ubjAI  (j1  j)1  jF1  jc1  j�1  j�1  j�1  j�1  j�1  j2  j.2  jK2  jh2  j�2  j�2  j�2  j�2  j�2  j3  j33  jP3  jm3  j�3  j�3  j�3  j�3  j�3  j4  j84  jU4  jr4  j�4  j�4  j�4  j�4  j5  j 5  j=5  jZ5  jw5  j�5  j�5  j�5  j�5  j6  j%6  jB6  j_6  j|6  j�6  t�����}�(jFI  ]�(j1  j)1  jF1  jc1  j�1  j�1  j�1  j�1  j�1  j2  j.2  jK2  jh2  j�2  j�2  j�2  j�2  j�2  j3  j33  jP3  jm3  j�3  j�3  j�3  j�3  j�3  j4  j84  jU4  jr4  j�4  j�4  j�4  j�4  j5  j 5  j=5  jZ5  jw5  j�5  j�5  j�5  j�5  j6  j%6  jB6  j_6  j|6  j�6  ejHI  NjII  hhK ��h��R�(KK2��h!�B�        �?                      �?              �?      �?              �?      �?       @      �?      @      @              @       @      @      @      @      @      @      @       @      @      @      $@       @      @       @       @      @      @      �?      @      @      @      @      �?      �?              �?              �?      �?                              �?      �?�t�bjPI  jQI  hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j>I  �remove���R�hQ�_container1�j[I  �ube�_autotitlepos���title�j�7  )��}�(h@�hANhBh�hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  �normal�j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nub�_left_title�j�7  )��}�(h@�hANhBh�hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G        j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  jI  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nub�_right_title�j�7  )��}�(h@�hANhBh�hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  jI  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nub�titleOffsetTrans�j�  �patch�j0+  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  jH+  jE+  �jF+  j7  jG+  jH+  jI+  jI  jP+  (G?�      G?�      G?�      G?�      t�jR+  G        jS+  K N��jU+  K N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  G        ji+  G        jm+  G?�      jq+  G?�      ju+  G        jv+  jw+  jx+  G?�      ub�axison���	fmt_xdata�N�	fmt_ydata�N�	_navigate���_navigate_mode�N�_shared_axes�}�h�]�(h�h>es�_twinned_axes�Nube�artists�]��lines�]�jFI  ]��texts�]��images�]��legends�]��subfigs�]��suppressComposite�N�_layout_engine�N�_fig_callbacks�hZ)��}�(h]]��dpi_changed�ah`hbhc}�heK hfNhg��ub�_canvas_callbacks�hZ)��}�(h]]�(�resize_event��
draw_event��key_press_event��key_release_event��button_press_event��button_release_event��scroll_event��motion_notify_event��
pick_event��figure_enter_event��figure_leave_event��axes_enter_event��axes_leave_event��close_event�eh`hbhc}�(j�I  }�K �matplotlib.backend_bases��_key_handler���sj�I  }�Kj�I  sj�I  }�(Kj�I  �_mouse_handler���Kh�hG�pick���R�uj�I  }�Kj�I  sj�I  }�(Kj�I  Kh�hGj�I  ��R�uj�I  }�Kj�I  suheKhfNhg��(K KKKKKKK�ub�_mouse_key_ids�]�(K KKKKKKe�_button_pick_id�K�_scroll_pick_id�K�bbox_inches�j�  �dpi_scale_trans�hό_dpi�G@Y      j�*  hҌfigbbox�hҌtransFigure�hՌtransSubfigure�h�j�I  j0+  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  (G?�      G?�      G?�      G?�      t�jE+  �jF+  j�I  jG+  jJ  jI+  j�I  jP+  jJ  jR+  G        jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  K ji+  K jm+  Kjq+  Kju+  G        jv+  jw+  jx+  G?�      ub�_original_dpi�G@Y      �subplotpars�hD�SubplotParams���)��}�(j'7  G?�      j�7  G?�(�\)j�8  G?�������jKF  G?�(�\)�wspace�G?ə������hspace�G?ə�����ub�_axstack�hD�
_AxesStack���)��}�(hB}�(h>Kh�Ku�_counter�Kub�_axobservers�hZ)��}�(h]Nh`hbhc}��_axes_change_event�}�sheKhfNhg��ub�number�K�__mpl_version__��3.7.2�ubhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�hGh���R�hjNhkNhlNhmNhnhohphs]�]�����hx�h�j�  j�*  h�)��}�(h�}�h�K h�hRj�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubj�*  h7j�*  j�*  j�*  j�*  j�*  }�(h~�h��uj�*  Nj�*  Nj�*  h�j�*  h�)��}�(h�}�h�Kh�hRj�  hhK ��h��R�(KKK��h!�C �?IoN�?���`C!⿡�Wۦ@ڜ��H��?�t�bj�  hhK ��h��R�(KK��h!�C�?IoN�? �iK?�t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �      �      ��      ���t�bubj�*  j�  j�*  jl  j�*  h�j�*  jt  j�*  h�j�*  h�j�*  j�  j�*  �matplotlib.gridspec��SubplotSpec���)��}�(�	_gridspec�jVJ  �GridSpec���)��}�(j'7  Nj�7  Nj�8  NjKF  NjJ  NjJ  NhChG�_nrows�K�_ncols�K�_row_height_ratios�]�Ka�_col_width_ratios�]�Kaub�num1�K �_num2�K ubj +  Nj+  j+  )��}�(j+  j
+  j(+  K j)+  K j*+  Kj++  Kubj,+  ]�(�matplotlib.collections��PathCollection���)��}�(h@�hANhBh>hChGhIj�  )��}�(h�}�h�Kh�hRh�NubhJ�hK�hL�hMG?�      hNj�  hONhP�hQ�Train $R^2 = 0.885$�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�jjJ  �remove���R�hjNhkNhlNhmNhnNhphs]�]�����hx��_A�N�_norm��matplotlib.colors��	Normalize���)��}�(�_vmin�N�_vmax�N�_clip��j�7  NhchZ)��}�(h]]��changed�ah`hbhc}�j�J  }�sheKhfNhg��ubub�_id_norm�K �cmap�j�J  �LinearSegmentedColormap���)��}�(�
monochrome��h8�Greys��N�M �	_rgba_bad�jH+  �_rgba_under�N�
_rgba_over�N�_i_under�M �_i_over�M�_i_bad�M�_isinit���colorbar_extend���_segmentdata�}�(�red�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�green�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�blue�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�alpha�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?�t�bu�_gamma�G?�      ub�colorbar�NhchZ)��}�(h]]�j�J  ah`hbhc}�heK hfNhg��ub�_us_linestyles�]�K N��aj�6  ]�h0h!C        ���R�N��a�_us_lw�hhK ��h��R�(KK��h!�C333333�?�t�b�_linewidths�j�J  �_face_is_mapped���_edge_is_mapped���_mapped_colors�NjC+  jD+  jI+  hhK ��h��R�(KKK��h!�C �?�������?TTTTTT�?      �?�t�b�_facecolors�hhK ��h��R�(KKK��h!�C �?�������?TTTTTT�?      �?�t�bjF+  �face��_edgecolors��face��_antialiaseds�hhK ��h��R�(KK��h�b1�����R�(K�|�NNNJ����J����K t�b�C�t�bj7  G@      �_urls�]�NajZ+  Nj8  Kj[+  Njb+  N�_offsets��numpy.ma.core��_mareconstruct���(j�J  �MaskedArray���hK ���b�t�R�(KMK��h!�B�!  ޯuŢ��?��m��������?�$�޻ۿ6Ah"���?�	B��?K�C.���?��'�3-���i�`��?�@'���?� �����? �H�?��AU�@��d/�����Az4@@e�Շb�����w��? l�Cy;U?�Hc�pw�? �c�ޭ�W�$K�!�?�ڵM�罿��_��? ����n?���@�l9�*�?sgn����?�;sSu�?IJɧrB�?X\X��<�?8���Y�@@Aߓ���?�� ,�@`j�Lg���h�Ҧ�?��]�?��>�1�?�#Z�?��.�zB ��?��=4��?<����@@l�a�����S��v@��[+����L3�? }�f���?n��`�i�?P�y$���6�>�$�?��+��?�0�@�r�����?,�+��� @8P:ӿ�e^��`�?�ړ�p�Qh��@@��G�_�?~A��@P�U��� %�ߩ@ �f�/F�?�w���?P~��vmȿ��|����?�ǆ�Nǖ?rB!���?�����ĵ��Xd}0�?��E�ð?�n�Lq�?H��#�?I��uY�?th��3\ٿ�N��9��?h��p0vȿ9�J���?`��u\Ơ?틞�d��?@k�0&�?�P��*�? BM<ª�?�bf�?p�!6Aa�?��n=�@ ���¥?�y�ث�@ F_N�v�s9��Z��? 8?�{���ˮt���?x�D-f пf�,]oA�? ��{��r��%|@ �~����K���\+�?�q�Y���?"���@@��ɫ��p�S��?����:������</�? �[�L������Dv��? ]V&�+�?�hL���?(�:��ܿ�Iȷ;�?����A"οhp �,�? ��2�1��|aA�\��?�:A	n���)ᔒ'�@���'���hze��?����A���g.��?0��[�ο\�Q"җ�?`����?~%O�@�W�$��?3�W���?��'��m�?�W飩@ � �-��?�O֔$@��#Z4,�?/h�5��?�&Z�?c=m_z�? ����s?=��#"�?@
�������0^�? mGKࢪ�1/�+��?Ps��뵿�՜�E@ ��0����B4i���@�`ll�?XӮ}JS�?@�邜�?�ܻ�'f@ iH̑�?��T�f�?H�8�B5�?�,�!��?�e�&1�?w�:��?'�:��?��#�{��?��G��$�?�5�ܜ�?xH����?屄�֔@`	c]�g�?G{	���?�@��u��?�����a�?����E׿U3V@&��?1at���d>��?�K%�r��p���w�?`ؒ�t��E�x�iN�?���@�?xY�9�?��ڈ��?�-Nڐ��?���ɿ?�[i3us�?\]'���ֿ��NȢ�?�t���?�guB��? *J���?�/M��.@��r���?������@ Z�
���?����
 @ ����
�?Y�@@���6��mN�s$��?ڜ��H��?>S�ܺ��?�35ȭ��?|�w�h�?@xĎ�v��J�T����?�yo>Fҿh����?�{;��?���>
�?D��\�������@�Q��L�?B'�� �?�&q���?"(�R|H�?����?D+��H�?� Z�D�?2��Ta��?��c�@ӿ�x�&���? Y49_��?��'2'@ >�\x�~�޷�` @�_��-5�?$N��q�? ��nk@�?�=u���@ +]a�n���9l�?P,��o���$���?1�V�ɿ�7�>� @���}RǿS�(#I @ /R��P׿DU,F�a�? �D耤Q����".��?�p|�zؿ".Y���?�q���?�sR�?�?��؊����9�D�@ ��O$��?�ǇPy��?`�ӻ�]���8ҵ��?��q|����2����?�^!�{ټ?�7��a�?`#z��i�?ni�8#� @�-�g��?׉:��@ �xP��?��=�Rt�?���<N�ӿ�2����@��Г���G��h�@ ��5e̕�e�ޡ�d@�{�{z���A��~+�?���{�=ȿt�},t#�?`��^�οnH���,@ K�,0���'���:�?��m�RS��������?���1��¿��-;P��?�M��ݿ��\�&�?P�����?��/>�?���O�οv��1
@ w@��?��%�E�? ���r?�X%� ��? ��D�?�A9�W�?H�I���?#��I�?趓�%ϿMd��p�?�Έ���?��c��@�`�&Z����i��@ I�We%��u3xÄ�@��_�͕��@�����@�a��9��?�u��x@��83wȿ��},K@ ��},K�?Zl�J�E@ P��뤿�^07J�?��s��?�u�tڄ�?���b�ڿC>�Tz��?���x�jڿ.`s�+@(��e!:п[�)L���?��.w��?.4 ��B@@z�߈������2p��?@���?�?���pm@�s�Y����qX��?���ú�? 1��'&�?�������?�3��?�Kl\�����i¿?�?Ppe}b�?&4���V�? n.����?8H���@ }�AT�?$g�Ku�? ��q�����c�@0��VͿz�67�?�O��?�T
�?(��z�Կ����� @�}���?�W<�d�?�U4z���?(|�W[��?`�Mܾ~̿��b,�@_�-ƒ�?i �U���?��(P�������Y�?��+:�0�?[D�I�?@H�[d���Q��&�?���U4пH�3�; @��`�ſs�{u�@ [6����?�6~vnT�?@k�g�F�?����@�,�)'�?�1�?x��p���?a�. � @ �c-���ȯ�F��?����?��<�+d�?��L����0�@���MnӤ������B�?���B�>�?�]�r�@�<��'�?Ă�I���?���x��?Q�飩��?ŝ>�z�?���_��@@�Kq�?]w�y @ �ݼ\���l�:�j�?`��C}D�?������?X��U%O�?��t�U�?�h蠒�?J=�S���?����?k����r @�J=�j¿����ʯ @�4}��9��R�L��? ��Ks���O�^:���?�>�?]e�?$=x��o�?�`��e6��Q'���� @ In�"��l�A\�? ��F��?�9@�!b������
��?8;��^�?7��kQ�? ٬��ݥ�4��u@���F�ޑ�8�뉐�?���j������@��R �S����b�]�@`y�eU%�?B�L�8e�? @��2����-��?�Y�TP����o+@�E,h��Ŀ�簮�?�E۷G��?���}b�@  ���\�4�K���?�?���G��xWxY���?�����8����f�P�?���7��?����\@PL���Z�?�&IzD�@ Pٶ����h�͙���?��[Y&_��W/>K��?�#_s�C�?0_���@��_���?	��0��?Ȋ"�(�?�d�8]@�����?�x�3��?p�%�ּ�?0��!���?b�"И�{ U�v��?`�(��ݧ��������?���T�f��WRr+��?���`C!⿤��]�?�X�U��wT�a��? ��<�~�s�o9'��? :�1���?�I��?�ǁu���q\e���?�>!��i��!� �D�?	�%�?n(܍q@@�zD�Q���!A���?0��˿˾�&+ @��8�ƿ6F���? ���ݔ�ݾe�0~�?O�j�ٿ�n�Ѧ�?xu�'�6�? ��^��?�,�����ˁz�?��T�A�?هt�K��?�RbT�?:���S�?0�Rgſo�Fq�? ~V1�e?~*=���@���ɘ�?h��b�O@ Z����?v�)��@`(�^xs�?��j���?`��I�A�?�2�zLH�?���$ĿrG�%���?@���'��4��i��? gJU���?�`�\-�?�J�Y�Կ��GX�-�?��?��l�?�a}�ݝ�? 0��������o!���?��qoJ�?����F @ =��1��?kP�PS�?��+�+&п�
�#�q@ r�YH����oH�@����@�?���!�$ @��:b�����mӐ�@�S�R�?�Rx׷�?`s��?/�	n@���G?��	�� @@8��#��?���e���?�0p����3�3!��?�������L(E���?������J���e@�v|(@B���}��ޔ�?��^AQyҿ"��/��?@t�i#E��p>=���@ ��c���?ȟM�"��?@�l���?^�b���? Q��N����#�?��??R����?���~��?��%b>�?QDZ@�c���?l�)^}l�?cu{ÿwm�d��?�� ������v[��?Щ�{]����.����?�o��X��?@�Y闧�? 0+��?l
8����?|��uO��?$�w��=�?� �;Y�����=�'�?��5iR��ϴui�� @p�ʿ"��_l @����%��c�:(�?D���,Կ���~@�5��rC˿����G4�?��e>����"^��b�?����?>��K��?���]��?}}�8ą�?���kA��?����?���ڳ��?�j�?��?@�|:�h��O�����?L1�Q&�?l�d�!�? :GFtп�n%m��?�tC(i��?��[���? �k��aT���g,$x�?@i��a��z��Tf��?��Ke�?��8��?��O�>ӿ�q�q"�? �5iDi�?<W�H1@�����Qÿk�5�
��?��#���?,��RG�@��m.u�?,��7KT@����D�?�)����?�Tߗ˚���p<@�? J���Ϝ?�Q	��?���!�A�?(=�����?@�D�?�ǳ��^�? �y��]��>4Y�#�?b7�S��?�k��@ �k�ă?��/�� �? ���<��*-P�e�?H�0jƿ*Qz���? kW�¶v��[w�Ek@��*��>�(���?����{���ǁ�D@@�o����2���?`g�<c(��:XJK���?`q��8�ÿ��:���?H=�ǂ�Ŀ��B=��? T;��v�@%|b���?h�V��?R��B�@��ǧ��?eM0%a�?`�\�Yۣ�$~F�׿@�C-{�֬�MB�rT��?0��Ŀ$���@ yF+:��[lJ�U�@`A¶���Xb�@`t���е���kRp@P�s|.̿*3����?��03���?�l���?`���힤?!y�m�@H^����п���I���? ��nظ���!;@���q.�?�S���?��}/�?R�N�;��?G�uO������w�?��Vt��x��J�W@���h����=�J�@@i����hf��>O�?���2 '�?^*�[�?x��o=H�?] {����?��qMg�?���w�4@�v�H��?1��z!}�?�!����?��|",� @ w�>��Ϳ��2�@�2�������!�=�?�I�AZ���A�A��@�Y�N�뮿����@��? L/Խ?%�&�@�X��(�?V	D�TF@ #�V!�?r��U�?P
��(��?+��O��?��f�?��?)4��g�? {�t�Q�?Hv6][��?���_}�����v��i�? �iK?��F���?���7R�?�Q����@�����?�n���@ �x0��?LRt�,��?�9�o����cx۳��?��Y��/�����s���? k�:���?�������?��7t=$�?�/����?�K�C��?�=$ny�@@$�i�ƿxMiA���?�kJe�?j(,=��?��p`�ò��4M����?��i��E�?z߅��?�Eu޽�(V��s��?`�f��-Ϳ���8ʦ�?@�HK��������\�?@
gj�ɪ���,�Z�?T����.п��vi��?`+b�Ʀ?���ٔ @h�)��Կo>n �@�jRjC@�?����b@ {�w�a��1Y�ۂ��? c�w��?DU��V�?x������?K.:�v�@��3nw�?(:N���?�.>��˿�C��)�?�E� ޴�?��_���?�AZ�| �?h�Y�,�@�&��.��?������?�?F08���H�D�?�%^#ڽ?CANsv��?0�4g׾?�"v����?@(b����?W��X�?�E/��S�?vʇ���@ AR�E�?x���3@��-ÿ��U��R @ O=�nĿh��E�?@k��p,�?U׶�?�5k��?���R��@����ִ���Ǒ����?����ڿ%�S���@����?z���P@ ���E����x��?�T~T�>ڿh���Hp�?8J�O�?���D�?�ê��&�?n��(�? ��bJaf�*��`�@@<��_��?�Y��^�?t����?���>D�?p���?��� ��?`�a�?<��(���?P-�i#ǿ��,�ݶ�?@�e<v�?DX�;�2@ �wm�{����ҏ@ Z��K���{���@�Z{8�S�?~>���@ ��kQm�����L�}�?Ȝ5�ſ���_��?�g&l���a}C��?�xWA�ț�-d��|�?����Ŀ��0�ێ�?@����?���$\�?�S���q��T�%��?�k8-v=���u}�e�?�[�p���?��@���Y���?qY@�q�? ��De?��b��@�|�y@JM�4@�?`����ѧ���tߴF�?HiXY�ſ$֠㩽�?�C��Sb��GP�uA��?�^��Ͳ?)8gL��?Rp��$�?�U�)�@��-���?��i�@��/�׿������? �I�cS��T,6t�@��AH�/���h�LHA@ �j�2*|?K��Q���? �e�Dx�ko_�C@�����
�?>��	dg�?���Jy^ο���I@ ���|M�?0��q@ ����=�����c��?��3�狿P�SY$R�? wBt�����d�?�=�a��?�`:��i�?P�,6�Ŀ*���-�?P�Twdn�? k����?�@F-:	̿�n����@ ������?��")���?��I��?��,��@@������?��(2��?`�	ſ~����?���ڞ��?�󚩭�@�^#��Q�?�"�,O�?p,2���?�P�(�@�E����?�~�NL�?�A,p%v���# �b�@�Ko�"?�?v��)�P�?�]�m�+�?`b#��@ &6R���?C|ޢC�? �I�op?���6�p�?�S\́�?�aP3�?�1��Ԍ��A�����?�=����¿ze� ��?�s��Hנ?���|H�?�$}͉��?��#����?�&-�[���'�o�? 
��a��ҕ,���?�S,tܦ?��^z7@�jy���¿g�L�־�?�l��H	ʿ;a1�[�?=���?���"1�?p�
$^�?Vz@��6�? �G����Ew��/�?��6bMԿ\���@ ��i�m?Ch��c��?`��q��?CW8�7d�?���'�wοNɹ-��?t8%�x�?j�p���?���\_K��B��j�@��:0��?���2���?��k�����p�O�E�?�	����ӿڄ�n�@�4J�[��?l�І @8c�xٿZjN��)�?�F&/�Lȿ�+C��?����ѿ7|����?��S�<��?��
���?���Jc��$�wP�&�?�P��?�����M@�:��5��?�4M@ G��^��%��?� �M
t��N���	@�p�ܽM�?3�e�@ �J��C�-���? ��l��r��Aɢ�@����?Zi�@���?`j��˦���2��?���9�í�������?@�Z�	w��6-:��?���T �?��,K�@@foeY��?���{���?��T��ÿ �Y�@ �Qg�_ƿ`�2���?0-�CQ�����Zs�?;�<���?1O�ν��?��^�ve�?�%pz�?���2����K��?@z>���DM6���?@$�2����Բ4��?�������?��ƅ��?�����5�����Mr�@��U�x��nޭ0���?p�n��^�?t:E4z�?�O��Ȱӿ̦�53w�?@c����Ϳ�����@ � !�����#f$��@��C�Щ��N�[t��?�%w���̿����@��A���п���G�? �q>P���^|$���? ~�ol��?;.I\m�?@�_�H��?+'�v� @`�$���?|z3V[
�? ,dN%���V!��@ �K�?�iJaP�?Ps��-��"-;�U@ q2��?"u7�k�?�(�E�Q��T�Zz�	@ ����s?�j��/ @�C�iaؿj��w�?��?��辿
��=I�?�Ba�@O�?�)��H$�?@3��i����s�2� @`���l��Uh�\�(�?`��aT꪿���%�? Rc�o&��4B���?��/"���B8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �Nt�b�_offset_transform�h�_paths�j&  )��}�(j)  hhK ��h��R�(KKK��h!�B�                �rSl��?      ࿉��e��?���֠ܿ�;f���?�;f��ֿ���֠�?���e�п      �?rSl���      �?              �?rSl��?���֠�?���e��?�;f���?�;f���?���e��?���֠�?rSl��?      �?              �?rSl���      �?���e�п���֠�?�;f��ֿ�;f���?���֠ܿ���e��?      �rSl��?      �              �rSl������֠ܿ���e�п�;f��ֿ�;f��ֿ���e�п���֠ܿrSl���      �              �              ࿔t�bj0  hhK ��h��R�(KK��h�u1�����R�(Kj�J  NNNJ����J����K t�b�CO�t�bj1  Kj2  G?�q�q��j3  �j4  �ub���_sizes�hhK ��h��R�(KK��h!�C     �H@�t�b�_transforms�hhK ��h��R�(KKKK��h!�CH�q�q#@                        �q�q#@                              �?�t�bubjmJ  )��}�(h@�hANhBh>hChGhIj�  )��}�(h�}�h�Kh�hRh�NubhJ�hK�hL�hMG?�      hNj   hONhP�hQ�Test $R^2 = 0.895$�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�jjJ  �remove���R�hjNhkNhlNhmNhnNhphs]�]�����hx�j�J  Nj�J  j�J  )��}�(j�J  Nj�J  Nj�J  �j�7  NhchZ)��}�(h]]�j�J  ah`hbhc}�j�J  }�sheKhfNhg��ububj�J  K j�J  j�J  )��}�(j�J  �h8j�J  j�J  M j�J  jH+  j�J  Nj�J  Nj�J  M j�J  Mj�J  Mj�J  �j�J  �j�J  j�J  j�J  G?�      ubj�J  NhchZ)��}�(h]]�j�J  ah`hbhc}�heK hfNhg��ubj�J  ]�K N��aj�6  ]�h0h!C        ���R�N��aj�J  hhK ��h��R�(KK��h!�C333333�?�t�bj�J  jSK  j�J  �j�J  �j�J  NjC+  jD+  jI+  hhK ��h��R�(KKK��h!�C �������?xxxxxx�?�������?      �?�t�bj�J  hhK ��h��R�(KKK��h!�C �������?xxxxxx�?�������?      �?�t�bjF+  �face�j�J  j�J  j�J  hhK ��h��R�(KK��j�J  �j�J  t�bj7  G@      j�J  ]�NajZ+  Nj8  Kj[+  Njb+  Nj�J  j�J  (j�J  hj�J  j�J  t�R�(KK�K��h!�B�  ���X6
�?���G��L�f�w�@ �m��?Ay���)@���I��?y����? J��z��?���2�@�Gх������~���?h��p� Ͽ\���h�@�u껌�?�?IoN�?��M:�/ڿ�����?@I�}?[ܚ���?�>I=��? ��-���? `|o���?35h�}�? �_�<V��m�a���? �A�e�W?�&�e-1�?@)�MSڙ���Wۦ@�&�G�:�?�,��%��?��qZ�/�?�yX?@ ����t¿`s�,FS�?`0Ϛ2�����+@ �WA+��L䣓B~�?@F,�Ò?8G��5@��~��/¿�0�֌@�?��I�f�?��	�#��?h[���F����0��?���C9t�?���) @ x���?��=���? �4Jn��.	
H��?pIP@��?O�j ��?��0�i��?>Hy��? |kȂ﾿������?����j�ѿ�
��9��?�޲�c�ÿ�~�-��?��`�#�?�}E���?�r�)��?��c�c� @kz�}տ��3sA��?������̿*\���k�?�m:0�̿�K6�v@ 9������:�Ӷ��? u`Jԑ?���t�@��E!��ſ�$49� �?�$�"]��а~�.R@ �7�"�?�׊��v�? }�8Jo�?��W��k�?��`��L�?.u_d��?Pn+��?�_�
�?�2��U��?��o���?P����?���l��@���Φ��?U�3Ĥ�@ "YF48��@�c��E�?�?>ҵӿT�3���@��Ԭ���?�J�F�@��}�]��$��Rsr�? )|����?vIP�7�? b<=,��?�����%@���ns�? M��&�? hj��4�?!�;�NJ�?���$Gǿ���YB@��Q�l���0;��N�?(Sk ���?n�>�?�a��?	ٸ�?�?X�һ��Ͽ�c�
 @\���ȿZ^Y3�@@6u��?��m�x�+�?���N�����"�,@@�fi��?E8ڡ� @�=,��ؿ�p�X@`*��ĪͿ��Z���? �X�v��K��e�i@ AP�e�?��`v҇�?`�Ll�ÿ�ޣ��? ���Y+�?�i��@ x�*p�?�Ő��@P�&J�ƿ9��@@�#�Q�?�!Z�[@ ]�� ���YQ�F�?���ɾ�W���N�?�{25v���������?��5�����)�����?Г���״���Ҧ|:�?�P�������~z@HM����? ���@��B{�8�?[d�I��?X��ÿ�������?�Ҍ:��п�J9+d�?�֘z��\'���@ ��nS��T�Z��? ���<z�?&0�+�-@ 8���?ta}��@�ot�i˦�zX�t�?�:��?S��,d%�? �-�k�7���/@�S�%�˲?2�㮅�?(k���?F�璣�@��唟��?����)��?�<�N��?`>�j��? 4���A��v��ψ@����f�?k��ȸ@ �1k�.�?�����5�?�44�����Z����? w��Œ�? �JEf @ i��̂��N%�<��?�t*��I�?��&�ʈ�?��S�?D��e'�?�~-J��M�_�$@ ��K�|�1.R����?P�Ca���R���? �N)Ȃ�?�=�M�?�w�nb�?vc�X]@�����?��{��?���U�?«#Ĕ��?P�mu��?�>��1��?0G��@���T�%@�y�%�ĿY�B��?H/Q�|(�?�D��@ d��-�?������@ V��0��?z��ϫ�@����YпLJ�����?��l��?0����s@���X���?� �:� @`Y��Rǿ�?����?��P6��?�կ��@��c� ���x��L�&�?@b���?���
��? a�I���?���	_�?`~��ɑ�?ƿ��I�@ �I�l�?q-EP�? \�~�1��@{M�	�? e���ʵ���Z,��?�Ōa�ѿ*yz`r�?(�R�J߿�H��I��?`Q=,��� �S�@�][$��?�Q��S@� �o�������@��j[2׿�UN����?@��-��?Gi�p�?��ѯV?����-^���?��%����B                                                                                                                                                                                                                                                                                  �Nt�bjK  h�jK  j&  )��}�(j)  hhK ��h��R�(KKK��h!�B�                �rSl��?      ࿉��e��?���֠ܿ�;f���?�;f��ֿ���֠�?���e�п      �?rSl���      �?              �?rSl��?���֠�?���e��?�;f���?�;f���?���e��?���֠�?rSl��?      �?              �?rSl���      �?���e�п���֠�?�;f��ֿ�;f���?���֠ܿ���e��?      �rSl��?      �              �rSl������֠ܿ���e�п�;f��ֿ�;f��ֿ���e�п���֠ܿrSl���      �              �              ࿔t�bj0  jK  j1  Kj2  G?�q�q��j3  �j4  �ub��jK  hhK ��h��R�(KK��h!�C     �H@�t�bj"K  hhK ��h��R�(KKKK��h!�CH�q�q#@                        �q�q#@                              �?�t�bubj�6  )��}�(h@�hANhBh>hChGhIj�  hJ�hK�hL�hMNhNj^  hONhP�hQ�_child2�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�jjJ  �remove���R�hjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j�6  j�6  j�6  )��}�(j�6  h�j�K  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  j�6  j#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  �j7  Kj7  K j7  ]�(K Kej7  ]�(K K ej�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�bj7  hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  j�  j5  j�  j7  �j7  Nubej7  ]�j!7  j$7  )��}�(j'7  j)7  )��}�(h@�hANhBh>hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  j'7  j=7  jk7  j8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C         ����p�        �J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububj�8  j)7  )��}�(h@�hANhBh>hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  j�8  j=7  jk7  j8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?����p�      �?�J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububj�7  j)7  )��}�(h@�hANhBh>hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  j�7  j=7  j�E  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jL7  �jM7  �jN7  jP7  )��}�(j'+  jU7  )��}�(jX7  h7jY7  �jZ7  Nj[7  Kj\7  hhK ��h��R�(KK��h!�C(      �?       @      @      @      $@�t�bjc7  hhK ��h��R�(KK
��h!�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�bjj7  �j=7  j�K  ubj}7  j�>  )��}�(j�>  Kj�>  K j�>  �j�7  �j�>  �j�>  K j�>  �%1.2f�j�>  �j�>  j�>  j�>  �j=7  j�K  j�7  hhK ��h��R�(KK
��h!�CP      �?      �?      �?      �?      �?      �?       @      @      @      @�t�bubj�7  �j�7  �ubjv7  jP7  )��}�(j'+  jz7  )��}�j=7  j�K  sbj}7  j7  )��}�(j=7  j�K  j�7  hhK ��h��R�(KK ��h!�j�6  t�bubj�7  �j�7  �ubhchZ)��}�(h]]�j�7  ah`hbhc}�j�7  }�K j�7  h�h>j�7  ��R���R�(j&L  h~��}�j�7  j�7  )��sNt�bssheKhfNhg��(K �ubj�7  �j�7  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  h0h!C      8@���R�j�7  �Predicted Value�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@&      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�7  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  h0h!C9��8�c9@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�7  G@      j7  Kj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  j�7  j�7  j�7  j�7  j�7  )��j�7  Nj�7  Nj 8  �j8  G?�      j8  ]�(jaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNjR  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�joL  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j`L  ��j7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�L  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j`L  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�L  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j`L  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j`L  j�  K j�7  �0.50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j`L  j�  Kj�7  j�L  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�L  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�L  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j3M  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�L  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�jOM  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j�L  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  j'  j5  j   j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�L  j�  K j�7  �0.75�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�L  j�  Kj�7  juM  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�M  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�M  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j�M  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  j>  j5  j;  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�M  j�  K j�7  �1.00�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�M  j�  Kj�7  j-N  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  jJN  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  ���      j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  jJN  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  jJN  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  jM  j5  jJ  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jJN  j�  K j�7  �1.25�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jJN  j�  Kj�7  j�N  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  jO  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  jO  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  jO  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  j\  j5  jY  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jO  j�  K j�7  �1.50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jO  j�  Kj�7  j�O  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�O  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�O  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j�O  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  jk  j5  jh  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�O  j�  K j�7  �1.75�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�O  j�  Kj�7  jUP  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C       @���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  jrP  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C       @�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C       @        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       @        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  jrP  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  jrP  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C       @       @�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C        @               @      �?�t�bj#  jz  j5  jw  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jrP  j�  K j�7  �2.00�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jrP  j�  Kj�7  jQ  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      @���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j*Q  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      @�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      @        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      @        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j*Q  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j*Q  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      @      @�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       @              @      �?�t�bj#  j�  j5  j�  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j*Q  j�  K j�7  �2.25�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j*Q  j�  Kj�7  j�Q  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      @���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�Q  ��j7  ]�K aj7  �j�  hhK ��h��R�(KK��h!�C      @�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      @        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      @        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�Q  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j�Q  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK��h!�C      @      @�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       @              @      �?�t�bj#  j�  j5  j�  j7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�Q  j�  K j�7  �2.50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�Q  j�  Kj�7  j}R  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubjaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      @���R�j8  �j�7  G        jm+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  jmL  jU+  jnL  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�R  ��j7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  G@ z�G�j7  Kj7  K j7  j�R  ��j7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  j�L  jU+  j�L  jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  j�R  ��j7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�R  j�  K j�7  �2.75�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�R  j�  Kj�7  jS  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@      ubejD>  ]�jaF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNjf  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        jm+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jIS  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�K aj7  ]�K aj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  NubjA8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j(8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jeS  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G        jY+  �j�6  j�7  j�6  G?�      j�6  j 7  j7  j7  j8  Kj7  Kj7  K j7  ]�K aj7  ]�Kaj7  �j�  Nj�  Nj7  Nj#  Nj5  Nj7  �j7  Nubj_8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  ja+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jR+  G?�      jS+  K N��jU+  G        N��jW+  j�6  j�6  �j�6  j67  j�6  j�6  )��}�(j�6  h�j�S  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njb+  j�6  j[+  ja+  j�6  �ubj�6  Nj�6  Nj�6  G@      jY+  �j�6  j�6  j�6  G        j�6  j 7  j7  j7  j7  Kj7  K j7  ]�(K K ej7  ]�(K Kej7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj7  �j7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jKF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  Kj�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�8  j�8  j�8  G@333333ubaj�H  j�7  ubj8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C �Ԓ.�p�?        �[8^@        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�NububjKF  j)7  )��}�(h@�hANhBh>hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  j57  jE+  �jF+  j67  jG+  j57  jI+  j7  jP+  jH+  jR+  G?�      jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  j;7  jb+  jg+  j<7  jKF  j=7  j�K  j8  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C �Ԓ.�p�?      �?�[8^@      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�NubububjI  j�K  jI  jk7  jP+  jI  jI  �jI  �jI  NjI  �hchZ)��}�(h]]�(jI  jI  jI  eh`hbhc}�heK hfNhg��ubjI  G?�������jI  G?�������jI  NjI  �j I  j#I  )��}�(j&I  h>j'I  j(I  ubj)I  j#I  )��}�(j&I  h>j'I  j,I  ubj-I  �j.I  j0I  )��}�j3I  j6I  )R�sbj8I  ]�j:I  Nj;I  h=}���j<I  �matplotlib.legend��Legend���)��}�(h@�hANhBh>hChGhIj�  )��}�(h�}�h�Kh�hRh�NubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�h>�_remove_legend���R�hjNhkNhlNhmNhnhohphs]�]�����hx��prop�j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ub�	_fontsize�G@$      j�I  ]�(j�7  )��}�(h@�hANhBh>hChGhIh��CompositeAffine2D���)��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}������j	T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?-؂-��{@                      �?�t�bubh�h�)��}�(h�}������j	T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?-؂-��{@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  jsJ  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�7  )��}�(h@�hANhBh>hChGhIjT  )��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}��Ы��j1T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?"""""Rz@                      �?�t�bubh�h�)��}�(h�}��Ы��j1T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?"""""Rz@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  j.K  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nube�legend_handles�]�(j0+  )��}�(h@�hANhBh>hChGhIjT  )��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}��Pq�j[T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH��8��8�?                        ��8��8�?                              �?�t�bubh�h�)��}�(h�}��Pq�j[T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        \����y@              �?-؂-��{@                      �?�t�bubh�hhK ��h��R�(KKK��h!�CH��8��8�?        \����y@        ��8��8�?-؂-��{@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQjsJ  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  (G?�G?ܜ�����G?�TTTTTTKt�jE+  �jF+  j�J  jG+  jT  jI+  j�J  jP+  jT  jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  G�       ji+  G�       jm+  G@4      jq+  G@      ju+  G        jv+  jw+  jx+  G?�      ubj0+  )��}�(h@�hANhBh>hChGhIjT  )��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}������j�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH��8��8�?                        ��8��8�?                              �?�t�bubh�h�)��}�(h�}������j�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        \����y@              �?"""""Rz@                      �?�t�bubh�hhK ��h��R�(KKK��h!�CH��8��8�?        \����y@        ��8��8�?"""""Rz@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQj.K  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  (G?�������G?�xxxxxxG?�������Kt�jE+  �jF+  �g�jG+  j�T  jI+  j�T  jP+  j�T  jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  G�       ji+  G�       jm+  G@4      jq+  G@      ju+  G        jv+  jw+  jx+  G?�      ube�_legend_title_box��matplotlib.offsetbox��TextArea���)��}�(j�7  j�7  )��}�(h@�hANhBh>hChGhIjT  )��}�(h�Kh�Kh�}�h�Kh�hRh�Nh�h�)��}�(h�}������j�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}������j�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�NubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubh@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�j�T  a�_offset�K K ���offset_transform�j�T  �_baseline_transform�j�T  �_multilinebaseline��ub�_custom_handler_map�N�	numpoints�K�markerscale�G?�      �scatterpoints�K�	borderpad�G?ٙ������labelspacing�G?�      �handlelength�G@       �handleheight�G?�ffffff�handletextpad�G?陙�����borderaxespad�G?�      �columnspacing�G@       �shadow��jaJ  K�_scatteryoffsets�hhK ��h��R�(KK��h!�C      �?�t�b�_legend_box�j�T  �VPacker���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�(j�T  j�T  �HPacker���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�j�T  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�(jU  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�(j�T  �DrawingArea���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�jYT  aj�T  h0h!C\����y@���R�h0h!C-؂-��{@���R����width�G@4      �height�G@      �xdescent�G        �ydescent�G        �_clip_children��j�T  jgT  �dpi_transform�j^T  ubj�T  )��}�(j�7  jT  h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�jT  aj�T  h0h!C@�~&f|@���R�h0h!C-؂-��{@���R���j�T  jT  j�T  jT  j�T  �ubej�T  h0h!C\����y@���R�h0h!C-؂-��{@���R���jAU  Nj@U  N�sep�G@       �pad�K �mode��fixed��align�j�7  ubjU  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�(j,U  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�j�T  aj�T  h0h!C\����y@���R�h0h!C"""""Rz@���R���j@U  G@4      jAU  G@      jBU  G        jCU  G        jDU  �j�T  j�T  jEU  j�T  ubj�T  )��}�(j�7  j/T  h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j,+  ]�j/T  aj�T  h0h!C@�~&f|@���R�h0h!C"""""Rz@���R���j�T  j4T  j�T  j=T  j�T  �ubej�T  h0h!C\����y@���R�h0h!C"""""Rz@���R���jAU  Nj@U  Nj`U  G@       jaU  K jbU  jcU  jdU  j�7  ubej�T  h0h!C\����y@���R�h0h!C-؂-��{@���R���jAU  Nj@U  Nj`U  G@      jaU  K jbU  jcU  jdU  j�7  ubaj�T  h0h!C\����y@���R�h0h!C-؂-��{@���R���jAU  Nj@U  Nj`U  G@4      jaU  K jbU  jcU  jdU  j�7  ubej�T  h�j�S  �_findoffset���R�jAU  Nj@U  Nj`U  G@      jaU  G@      jbU  jcU  jdU  j�7  ub�isaxes���parent�h>�_loc_used_default���_outside_loc�N�_mode�N�_bbox_to_anchor�N�legendPatch�j.+  �FancyBboxPatch���)��}�(h@�hANhBh>hChGhIj�S  hJ�hK�hL�hMG?陙����hNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhl�hmNhnhohphs]�]�����hx�jC+  (G?陙����G?陙����G?陙����G?陙����t�jE+  �jF+  �0.8�jG+  j�U  jI+  jI  jP+  (G?�      G?�      G?�      G?陙����t�jR+  G?�333333jS+  K N��jU+  G        N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  j�  h0h!C���
�y@���R�j�  h0h!C�>�>�y@���R�jm+  h0h!C���c@���R�jq+  h0h!C�`��K@���R��_bbox_transmuter�j.+  �BoxStyle.Round���)��}�(jaU  G        �rounding_size�G?ə�����ub�_mutation_scale�G@+�q�r�_mutation_aspect�Kub�
_alignment�j�7  �_legend_handle_box�jU  �	_loc_real�K �
_draggable�Nubj=I  ]�jpI  �jqI  j�7  )��}�(h@�hANhBh>hChGhIjH  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  �$Residuals for LinearRegression Model�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  jI  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  �center�j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�I  j�7  )��}�(h@�hANhBh>hChGhIjN  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G        j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  jI  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j'7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�I  j�7  )��}�(h@�hANhBh>hChGhIjQ  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  jI  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  Nubj�I  jK  j�I  j0+  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jC+  jH+  jE+  �jF+  j7  jG+  jH+  jI+  jI  jP+  j�I  jR+  G        jS+  K N��jU+  K N��jW+  jX+  jY+  �jZ+  Nj[+  ja+  jb+  jg+  jh+  G        ji+  G        jm+  G?�      jq+  G?�      ju+  G        jv+  jw+  jx+  G?�      ubj�I  �j�I  Nj�I  Nj�I  �j�I  Nj�I  }�h�]�(h�h>esj�I  Nubj+  Nj�7  N�color�NjqI  N�colors�}�(�train_point�j�J  �
test_point�j�T  j�E  j�6  u�hist���qqplot���_hax�h��_labels�]�(jsJ  j.K  e�_colors�]�(j�J  j�T  e�alphas�}�(jV  G?�      jV  G?�      u�train_score_�h0h!Cglk�T�?���R��test_score_�h0h!C�W�ע�?���R�ub.